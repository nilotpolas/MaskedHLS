module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    r6,
    r7,
    r8,
    r9,
    r10,
    r11,
    r12,
    r13,
    r14,
    r15,
    r16,
    r17,
    r18,
    r19,
    r20,
    r21,
    r22,
    r23,
    r24,
    r25,
    r26,
    r27,
    r28,
    r29,
    r30,
    r31,
    r32,
    r33,
    r34,
    r35,
    r36,
    r37,
    r38,
    r39,
    r40,
    r41,
    r42,
    r43,
    r44,
    r45,
    r46,
    r47,
    r48,
    r49,
    r50,
    r51,
    r52,
    r53,
    r54,
    r55,
    r56,
    r57,
    r58,
    r59,
    r60,
    r61,
    r62,
    r63,
    r64,
    r65,
    r66,
    r67,
    r68,
    r69,
    r70,
    r71,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1
);
//input [7:0]S
    input clk;
    input [7:0]  t0;
    input [7:0]  t1;
    input [7:0]  r0;
    input [7:0]  r1;
    input [7:0]  r2;
    input [7:0]  r3;
    input [7:0]  r4;
    input [7:0]  r5;
    input [7:0]  r6;
    input [7:0]  r7;
    input [7:0]  r8;
    input [7:0]  r9;
    input [7:0]  r10;
    input [7:0]  r11;
    input [7:0]  r12;
    input [7:0]  r13;
    input [7:0]  r14;
    input [7:0]  r15;
    input [7:0]  r16;
    input [7:0]  r17;
    input [7:0]  r18;
    input [7:0]  r19;
    input [7:0]  r20;
    input [7:0]  r21;
    input [7:0]  r22;
    input [7:0]  r23;
    input [7:0]  r24;
    input [7:0]  r25;
    input [7:0]  r26;
    input [7:0]  r27;
    input [7:0]  r28;
    input [7:0]  r29;
    input [7:0]  r30;
    input [7:0]  r31;
    input [7:0]  r32;
    input [7:0]  r33;
    input [7:0]  r34;
    input [7:0]  r35;
    input [7:0]  r36;
    input [7:0]  r37;
    input [7:0]  r38;
    input [7:0]  r39;
    input [7:0]  r40;
    input [7:0]  r41;
    input [7:0]  r42;
    input [7:0]  r43;
    input [7:0]  r44;
    input [7:0]  r45;
    input [7:0]  r46;
    input [7:0]  r47;
    input [7:0]  r48;
    input [7:0]  r49;
    input [7:0]  r50;
    input [7:0]  r51;
    input [7:0]  r52;
    input [7:0]  r53;
    input [7:0]  r54;
    input [7:0]  r55;
    input [7:0]  r56;
    input [7:0]  r57;
    input [7:0]  r58;
    input [7:0]  r59;
    input [7:0]  r60;
    input [7:0]  r61;
    input [7:0]  r62;
    input [7:0]  r63;
    input [7:0]  r64;
    input [7:0]  r65;
    input [7:0]  r66;
    input [7:0]  r67;
    input [7:0]  r68;
    input [7:0]  r69;
    input [7:0]  r70;
    input [7:0]  r71;
    input [7:0]  dec_0;
    input [7:0]  dec_1;
    input [7:0]  dec_255;
    input [7:0]  dec_169;
    input [7:0]  dec_129;
    input [7:0]  dec_9;
    input [7:0]  dec_72;
    input [7:0]  dec_242;
    input [7:0]  dec_243;
    input [7:0]  dec_152;
    input [7:0]  dec_240;
    input [7:0]  dec_4;
    input [7:0]  dec_15;
    input [7:0]  dec_12;
    input [7:0]  dec_2;
    input [7:0]  dec_3;
    input [7:0]  dec_16;
    input [7:0]  dec_36;
    input [7:0]  dec_220;
    input [7:0]  dec_11;
    input [7:0]  dec_158;
    input [7:0]  dec_45;
    input [7:0]  dec_88;
    input [7:0]  dec_99;
//OUTPUTS
    output reg [7:0]  y0;
    output reg [7:0]  y1;
//Intermediate values
    wire [7:0] dec_99_inp;
    wire [7:0] dec_88_inp;
    wire [7:0] dec_45_inp;
    wire [7:0] dec_158_inp;
    wire [7:0] dec_11_inp;
    wire [7:0] dec_220_inp;
    wire [7:0] dec_36_inp;
    wire [7:0] dec_16_inp;
    wire [7:0] dec_3_inp;
    wire [7:0] dec_2_inp;
    wire [7:0] dec_12_inp;
    wire [7:0] dec_15_inp;
    wire [7:0] dec_4_inp;
    wire [7:0] dec_240_inp;
    wire [7:0] dec_152_inp;
    wire [7:0] dec_243_inp;
    wire [7:0] dec_242_inp;
    wire [7:0] dec_72_inp;
    wire [7:0] dec_9_inp;
    wire [7:0] dec_129_inp;
    wire [7:0] dec_169_inp;
    wire [7:0] dec_255_inp;
    wire [7:0] dec_1_inp;
    wire [7:0] dec_0_inp;
    wire [7:0] t0_inp;
    wire [7:0] t1_inp;
    wire [7:0] r0_inp;
    wire [7:0] r1_inp;
    wire [7:0] r2_inp;
    wire [7:0] r3_inp;
    wire [7:0] r4_inp;
    wire [7:0] r5_inp;
    wire [7:0] r6_inp;
    wire [7:0] r7_inp;
    wire [7:0] r8_inp;
    wire [7:0] r9_inp;
    wire [7:0] r10_inp;
    wire [7:0] r11_inp;
    wire [7:0] r12_inp;
    wire [7:0] r13_inp;
    wire [7:0] r14_inp;
    wire [7:0] r15_inp;
    wire [7:0] r16_inp;
    wire [7:0] r17_inp;
    wire [7:0] r18_inp;
    wire [7:0] r19_inp;
    wire [7:0] r20_inp;
    wire [7:0] r21_inp;
    wire [7:0] r22_inp;
    wire [7:0] r23_inp;
    wire [7:0] r24_inp;
    wire [7:0] r25_inp;
    wire [7:0] r26_inp;
    wire [7:0] r27_inp;
    wire [7:0] r28_inp;
    wire [7:0] r29_inp;
    wire [7:0] r30_inp;
    wire [7:0] r31_inp;
    wire [7:0] r32_inp;
    wire [7:0] r33_inp;
    wire [7:0] r34_inp;
    wire [7:0] r35_inp;
    wire [7:0] r36_inp;
    wire [7:0] r37_inp;
    wire [7:0] r38_inp;
    wire [7:0] r39_inp;
    wire [7:0] r40_inp;
    wire [7:0] r41_inp;
    wire [7:0] r42_inp;
    wire [7:0] r43_inp;
    wire [7:0] r44_inp;
    wire [7:0] r45_inp;
    wire [7:0] r46_inp;
    wire [7:0] r47_inp;
    wire [7:0] r48_inp;
    wire [7:0] r49_inp;
    wire [7:0] r50_inp;
    wire [7:0] r51_inp;
    wire [7:0] r52_inp;
    wire [7:0] r53_inp;
    wire [7:0] r54_inp;
    wire [7:0] r55_inp;
    wire [7:0] r56_inp;
    wire [7:0] r57_inp;
    wire [7:0] r58_inp;
    wire [7:0] r59_inp;
    wire [7:0] r60_inp;
    wire [7:0] r61_inp;
    wire [7:0] r62_inp;
    wire [7:0] r63_inp;
    wire [7:0] r64_inp;
    wire [7:0] r65_inp;
    wire [7:0] r66_inp;
    wire [7:0] r67_inp;
    wire [7:0] r68_inp;
    wire [7:0] r69_inp;
    wire [7:0] r70_inp;
    wire [7:0] r71_inp;
    wire [7:0] y_G256_newbasis0;
    wire [7:0] tempy1_G256_newbasis0;
    wire [7:0] cond1_G256_newbasis0;
    wire [7:0] negCond1_G256_newbasis0;
    wire [7:0] yxorb1_G256_newbasis0;
    wire [7:0] ny1_G256_newbasis0;
    wire [7:0] tempyIntoNegCond1_G256_newbasis0;
    wire [7:0] y1_G256_newbasis0;
    wire [7:0] x1_G256_newbasis0;
    wire [7:0] tempy2_G256_newbasis0;
    wire [7:0] cond2_G256_newbasis0;
    wire [7:0] negCond2_G256_newbasis0;
    wire [7:0] yxorb2_G256_newbasis0;
    wire [7:0] ny2_G256_newbasis0;
    wire [7:0] tempyIntoNegCond2_G256_newbasis0;
    wire [7:0] y2_G256_newbasis0;
    wire [7:0] x2_G256_newbasis0;
    wire [7:0] tempy3_G256_newbasis0;
    wire [7:0] cond3_G256_newbasis0;
    wire [7:0] negCond3_G256_newbasis0;
    wire [7:0] yxorb3_G256_newbasis0;
    wire [7:0] ny3_G256_newbasis0;
    wire [7:0] tempyIntoNegCond3_G256_newbasis0;
    wire [7:0] y3_G256_newbasis0;
    wire [7:0] x3_G256_newbasis0;
    wire [7:0] tempy4_G256_newbasis0;
    wire [7:0] cond4_G256_newbasis0;
    wire [7:0] negCond4_G256_newbasis0;
    wire [7:0] yxorb4_G256_newbasis0;
    wire [7:0] ny4_G256_newbasis0;
    wire [7:0] tempyIntoNegCond4_G256_newbasis0;
    wire [7:0] y4_G256_newbasis0;
    wire [7:0] x4_G256_newbasis0;
    wire [7:0] tempy5_G256_newbasis0;
    wire [7:0] cond5_G256_newbasis0;
    wire [7:0] negCond5_G256_newbasis0;
    wire [7:0] yxorb5_G256_newbasis0;
    wire [7:0] ny5_G256_newbasis0;
    wire [7:0] tempyIntoNegCond5_G256_newbasis0;
    wire [7:0] y5_G256_newbasis0;
    wire [7:0] x5_G256_newbasis0;
    wire [7:0] tempy6_G256_newbasis0;
    wire [7:0] cond6_G256_newbasis0;
    wire [7:0] negCond6_G256_newbasis0;
    wire [7:0] yxorb6_G256_newbasis0;
    wire [7:0] ny6_G256_newbasis0;
    wire [7:0] tempyIntoNegCond6_G256_newbasis0;
    wire [7:0] y6_G256_newbasis0;
    wire [7:0] x6_G256_newbasis0;
    wire [7:0] tempy7_G256_newbasis0;
    wire [7:0] cond7_G256_newbasis0;
    wire [7:0] negCond7_G256_newbasis0;
    wire [7:0] yxorb7_G256_newbasis0;
    wire [7:0] ny7_G256_newbasis0;
    wire [7:0] tempyIntoNegCond7_G256_newbasis0;
    wire [7:0] y7_G256_newbasis0;
    wire [7:0] x7_G256_newbasis0;
    wire [7:0] tempy8_G256_newbasis0;
    wire [7:0] cond8_G256_newbasis0;
    wire [7:0] negCond8_G256_newbasis0;
    wire [7:0] yxorb8_G256_newbasis0;
    wire [7:0] ny8_G256_newbasis0;
    wire [7:0] tempyIntoNegCond8_G256_newbasis0;
    wire [7:0] y8_G256_newbasis0;
    wire [7:0] z3225_assgn3225;
    reg [7:0] z3225_assgn32250;
    reg [7:0] z3225_assgn32251;
    reg [7:0] z3225_assgn32252;
    reg [7:0] z3225_assgn32253;
    reg [7:0] z3225_assgn32254;
    reg [7:0] x8_G256_newbasis0;
    wire [7:0] t2;
    wire [7:0] z_y_G256_newbasis0;
    wire [7:0] z_tempy1_G256_newbasis0;
    wire [7:0] z_cond1_G256_newbasis0;
    wire [7:0] z_negCond1_G256_newbasis0;
    wire [7:0] z_yxorb1_G256_newbasis0;
    wire [7:0] z_ny1_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond1_G256_newbasis0;
    wire [7:0] z_y1_G256_newbasis0;
    wire [7:0] z_x1_G256_newbasis0;
    wire [7:0] z_tempy2_G256_newbasis0;
    wire [7:0] z_cond2_G256_newbasis0;
    wire [7:0] z_negCond2_G256_newbasis0;
    wire [7:0] z_yxorb2_G256_newbasis0;
    wire [7:0] z_ny2_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond2_G256_newbasis0;
    wire [7:0] z_y2_G256_newbasis0;
    wire [7:0] z_x2_G256_newbasis0;
    wire [7:0] z_tempy3_G256_newbasis0;
    wire [7:0] z_cond3_G256_newbasis0;
    wire [7:0] z_negCond3_G256_newbasis0;
    wire [7:0] z_yxorb3_G256_newbasis0;
    wire [7:0] z_ny3_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond3_G256_newbasis0;
    wire [7:0] z_y3_G256_newbasis0;
    wire [7:0] z_x3_G256_newbasis0;
    wire [7:0] z_tempy4_G256_newbasis0;
    wire [7:0] z_cond4_G256_newbasis0;
    wire [7:0] z_negCond4_G256_newbasis0;
    wire [7:0] z_yxorb4_G256_newbasis0;
    wire [7:0] z_ny4_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond4_G256_newbasis0;
    wire [7:0] z_y4_G256_newbasis0;
    wire [7:0] z_x4_G256_newbasis0;
    wire [7:0] z_tempy5_G256_newbasis0;
    wire [7:0] z_cond5_G256_newbasis0;
    wire [7:0] z_negCond5_G256_newbasis0;
    wire [7:0] z_yxorb5_G256_newbasis0;
    wire [7:0] z_ny5_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond5_G256_newbasis0;
    wire [7:0] z_y5_G256_newbasis0;
    wire [7:0] z_x5_G256_newbasis0;
    wire [7:0] z_tempy6_G256_newbasis0;
    wire [7:0] z_cond6_G256_newbasis0;
    wire [7:0] z_negCond6_G256_newbasis0;
    wire [7:0] z_yxorb6_G256_newbasis0;
    wire [7:0] z_ny6_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond6_G256_newbasis0;
    wire [7:0] z_y6_G256_newbasis0;
    wire [7:0] z_x6_G256_newbasis0;
    wire [7:0] z_tempy7_G256_newbasis0;
    wire [7:0] z_cond7_G256_newbasis0;
    wire [7:0] z_negCond7_G256_newbasis0;
    wire [7:0] z_yxorb7_G256_newbasis0;
    wire [7:0] z_ny7_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond7_G256_newbasis0;
    wire [7:0] z_y7_G256_newbasis0;
    wire [7:0] z_x7_G256_newbasis0;
    wire [7:0] z_tempy8_G256_newbasis0;
    wire [7:0] z_cond8_G256_newbasis0;
    wire [7:0] z_negCond8_G256_newbasis0;
    wire [7:0] z_yxorb8_G256_newbasis0;
    wire [7:0] z_ny8_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond8_G256_newbasis0;
    wire [7:0] z_y8_G256_newbasis0;
    wire [7:0] z3357_assgn3357;
    reg [7:0] z3357_assgn33570;
    reg [7:0] z3357_assgn33571;
    reg [7:0] z3357_assgn33572;
    reg [7:0] z3357_assgn33573;
    reg [7:0] z3357_assgn33574;
    reg [7:0] z_x8_G256_newbasis0;
    wire [7:0] t3;
    wire [7:0] a0_0_G256_inv0;
    wire [7:0] a1_0_G256_inv0;
    wire [7:0] a0_G256_inv0;
    wire [7:0] a1_G256_inv0;
    wire [7:0] b0_G256_inv0;
    wire [7:0] b1_G256_inv0;
    wire [7:0] a0xorb0_G256_inv0;
    wire [7:0] a1xorb1_G256_inv0;
    wire [7:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] c0_G256_inv0;
    wire [7:0] c1_G256_inv0;
    wire [7:0] r00_G16_mul0_G256_inv0;
    wire [7:0] v_r1_G16_mul0_G256_inv0;
    wire [7:0] r20_G16_mul0_G256_inv0;
    wire [7:0] r30_G16_mul0_G256_inv0;
    wire [7:0] r40_G16_mul0_G256_inv0;
    wire [7:0] r50_G16_mul0_G256_inv0;
    wire [7:0] r60_G16_mul0_G256_inv0;
    wire [7:0] r70_G16_mul0_G256_inv0;
    wire [7:0] r80_G16_mul0_G256_inv0;
    wire [7:0] r90_G16_mul0_G256_inv0;
    wire [7:0] r100_G16_mul0_G256_inv0;
    wire [7:0] r110_G16_mul0_G256_inv0;
    wire [7:0] r120_G16_mul0_G256_inv0;
    wire [7:0] r130_G16_mul0_G256_inv0;
    wire [7:0] r140_G16_mul0_G256_inv0;
    wire [7:0] r150_G16_mul0_G256_inv0;
    wire [7:0] r160_G16_mul0_G256_inv0;
    wire [7:0] r170_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G16_mul0_G256_inv0;
    wire [7:0] a0_G16_mul0_G256_inv0;
    wire [7:0] a1_G16_mul0_G256_inv0;
    wire [7:0] b0_G16_mul0_G256_inv0;
    wire [7:0] b1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G16_mul0_G256_inv0;
    wire [7:0] c0_G16_mul0_G256_inv0;
    wire [7:0] c1_G16_mul0_G256_inv0;
    wire [7:0] d0_G16_mul0_G256_inv0;
    wire [7:0] d1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc10_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc10_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc10_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc11_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc11_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc11_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc11_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc12_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc12_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc12_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc12_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] z3661_assgn3661;
    reg [7:0] z3661_assgn36610;
    reg [7:0] z761_assgn761;
    wire [7:0] p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] z3665_assgn3665;
    reg [7:0] z3665_assgn36650;
    reg [7:0] z763_assgn763;
    wire [7:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G16_mul0_G256_inv0;
    wire [7:0] e1_G16_mul0_G256_inv0;
    wire [7:0] z3673_assgn3673;
    reg [7:0] z3673_assgn36730;
    reg [7:0] z769_assgn769;
    wire [7:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3677_assgn3677;
    reg [7:0] z3677_assgn36770;
    reg [7:0] z771_assgn771;
    wire [7:0] a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3681_assgn3681;
    reg [7:0] z3681_assgn36810;
    reg [7:0] z773_assgn773;
    wire [7:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3685_assgn3685;
    reg [7:0] z3685_assgn36850;
    reg [7:0] z775_assgn775;
    wire [7:0] a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3689_assgn3689;
    reg [7:0] z3689_assgn36890;
    reg [7:0] z777_assgn777;
    wire [7:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3693_assgn3693;
    reg [7:0] z3693_assgn36930;
    reg [7:0] z779_assgn779;
    wire [7:0] b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3705_assgn3705;
    reg [7:0] z3705_assgn37050;
    reg [7:0] z789_assgn789;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3709_assgn3709;
    reg [7:0] z3709_assgn37090;
    reg [7:0] z791_assgn791;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] e01_G16_mul0_G256_inv0;
    wire [7:0] e11_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc10_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc10_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc10_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc11_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc11_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc11_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc11_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc12_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc12_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc12_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc12_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] z3841_assgn3841;
    reg [7:0] z3841_assgn38410;
    reg [7:0] z921_assgn921;
    wire [7:0] p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] z3845_assgn3845;
    reg [7:0] z3845_assgn38450;
    reg [7:0] z923_assgn923;
    wire [7:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G16_mul0_G256_inv0;
    wire [7:0] p0_G16_mul0_G256_inv0;
    wire [7:0] p1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc10_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc10_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc10_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc11_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc11_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc11_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc11_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc12_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] r10_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] i1_hpc12_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_hpc12_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_hpc12_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] z3981_assgn3981;
    reg [7:0] z3981_assgn39810;
    reg [7:0] z1057_assgn1057;
    wire [7:0] p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] z3985_assgn3985;
    reg [7:0] z3985_assgn39850;
    reg [7:0] z1059_assgn1059;
    wire [7:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G16_mul0_G256_inv0;
    wire [7:0] q0_G16_mul0_G256_inv0;
    wire [7:0] q1_G16_mul0_G256_inv0;
    wire [7:0] z3997_assgn3997;
    reg [7:0] z3997_assgn39970;
    reg [7:0] z1069_assgn1069;
    wire [7:0] p0ls2_G16_mul0_G256_inv0;
    wire [7:0] z4001_assgn4001;
    reg [7:0] z4001_assgn40010;
    reg [7:0] z1071_assgn1071;
    wire [7:0] p1ls2_G16_mul0_G256_inv0;
    wire [7:0] d0_G256_inv0;
    wire [7:0] d1_G256_inv0;
    wire [7:0] z4009_assgn4009;
    reg [7:0] z4009_assgn40090;
    reg [7:0] z1078_assgn1078;
    wire [7:0] c0xord0_G256_inv0;
    wire [7:0] z4013_assgn4013;
    reg [7:0] z4013_assgn40130;
    reg [7:0] z1080_assgn1080;
    wire [7:0] c1xord1_G256_inv0;
    wire [7:0] r00_G16_inv0_G256_inv0;
    wire [7:0] v_r1_G16_inv0_G256_inv0;
    wire [7:0] r20_G16_inv0_G256_inv0;
    wire [7:0] r30_G16_inv0_G256_inv0;
    wire [7:0] r40_G16_inv0_G256_inv0;
    wire [7:0] r50_G16_inv0_G256_inv0;
    wire [7:0] r60_G16_inv0_G256_inv0;
    wire [7:0] r70_G16_inv0_G256_inv0;
    wire [7:0] r80_G16_inv0_G256_inv0;
    wire [7:0] r90_G16_inv0_G256_inv0;
    wire [7:0] r100_G16_inv0_G256_inv0;
    wire [7:0] r110_G16_inv0_G256_inv0;
    wire [7:0] r120_G16_inv0_G256_inv0;
    wire [7:0] r130_G16_inv0_G256_inv0;
    wire [7:0] r140_G16_inv0_G256_inv0;
    wire [7:0] r150_G16_inv0_G256_inv0;
    wire [7:0] r160_G16_inv0_G256_inv0;
    wire [7:0] r170_G16_inv0_G256_inv0;
    wire [7:0] z4053_assgn4053;
    reg [7:0] z4053_assgn40530;
    reg [7:0] z1117_assgn1117;
    wire [7:0] a0_0_G16_inv0_G256_inv0;
    wire [7:0] z4057_assgn4057;
    reg [7:0] z4057_assgn40570;
    reg [7:0] z1119_assgn1119;
    wire [7:0] a1_0_G16_inv0_G256_inv0;
    wire [7:0] z4061_assgn4061;
    reg [7:0] z4061_assgn40610;
    reg [7:0] z1121_assgn1121;
    wire [7:0] a0_G16_inv0_G256_inv0;
    wire [7:0] z4065_assgn4065;
    reg [7:0] z4065_assgn40650;
    reg [7:0] z1123_assgn1123;
    wire [7:0] a1_G16_inv0_G256_inv0;
    wire [7:0] z4069_assgn4069;
    reg [7:0] z4069_assgn40690;
    reg [7:0] z1125_assgn1125;
    wire [7:0] b0_G16_inv0_G256_inv0;
    wire [7:0] z4073_assgn4073;
    reg [7:0] z4073_assgn40730;
    reg [7:0] z1127_assgn1127;
    wire [7:0] b1_G16_inv0_G256_inv0;
    wire [7:0] a0xorb0_G16_inv0_G256_inv0;
    wire [7:0] a1xorb1_G16_inv0_G256_inv0;
    wire [7:0] z4081_assgn4081;
    reg [7:0] z4081_assgn40810;
    reg [7:0] z1133_assgn1133;
    wire [7:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4085_assgn4085;
    reg [7:0] z4085_assgn40850;
    reg [7:0] z1135_assgn1135;
    wire [7:0] a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4089_assgn4089;
    reg [7:0] z4089_assgn40890;
    reg [7:0] z1137_assgn1137;
    wire [7:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4093_assgn4093;
    reg [7:0] z4093_assgn40930;
    reg [7:0] z1139_assgn1139;
    wire [7:0] a1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4097_assgn4097;
    reg [7:0] z4097_assgn40970;
    reg [7:0] z1141_assgn1141;
    wire [7:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4101_assgn4101;
    reg [7:0] z4101_assgn41010;
    reg [7:0] z1143_assgn1143;
    wire [7:0] b1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4105_assgn4105;
    reg [7:0] z4105_assgn41050;
    reg [7:0] z1145_assgn1145;
    wire [7:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4109_assgn4109;
    reg [7:0] z4109_assgn41090;
    reg [7:0] z1147_assgn1147;
    wire [7:0] b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G16_inv0_G256_inv0;
    wire [7:0] z4117_assgn4117;
    reg [7:0] z4117_assgn41170;
    reg [7:0] z1153_assgn1153;
    wire [7:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4121_assgn4121;
    reg [7:0] z4121_assgn41210;
    reg [7:0] z1155_assgn1155;
    wire [7:0] a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4125_assgn4125;
    reg [7:0] z4125_assgn41250;
    reg [7:0] z1157_assgn1157;
    wire [7:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4129_assgn4129;
    reg [7:0] z4129_assgn41290;
    reg [7:0] z1159_assgn1159;
    wire [7:0] a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4133_assgn4133;
    reg [7:0] z4133_assgn41330;
    reg [7:0] z1161_assgn1161;
    wire [7:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4137_assgn4137;
    reg [7:0] z4137_assgn41370;
    reg [7:0] z1163_assgn1163;
    wire [7:0] b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4149_assgn4149;
    reg [7:0] z4149_assgn41490;
    reg [7:0] z1173_assgn1173;
    wire [7:0] p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4153_assgn4153;
    reg [7:0] z4153_assgn41530;
    reg [7:0] z1175_assgn1175;
    wire [7:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] c0_G16_inv0_G256_inv0;
    wire [7:0] c1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4173_assgn4173;
    reg [7:0] z4173_assgn41730;
    reg [7:0] z1193_assgn1193;
    wire [7:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4177_assgn4177;
    reg [7:0] z4177_assgn41770;
    reg [7:0] z1195_assgn1195;
    wire [7:0] a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4181_assgn4181;
    reg [7:0] z4181_assgn41810;
    reg [7:0] z1197_assgn1197;
    wire [7:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4185_assgn4185;
    reg [7:0] z4185_assgn41850;
    reg [7:0] z1199_assgn1199;
    wire [7:0] a1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4189_assgn4189;
    reg [7:0] z4189_assgn41890;
    reg [7:0] z1201_assgn1201;
    wire [7:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4193_assgn4193;
    reg [7:0] z4193_assgn41930;
    reg [7:0] z1203_assgn1203;
    wire [7:0] b1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4197_assgn4197;
    reg [7:0] z4197_assgn41970;
    reg [7:0] z1205_assgn1205;
    wire [7:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4201_assgn4201;
    reg [7:0] z4201_assgn42010;
    reg [7:0] z1207_assgn1207;
    wire [7:0] c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4205_assgn4205;
    reg [7:0] z4205_assgn42050;
    reg [7:0] z1209_assgn1209;
    wire [7:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4209_assgn4209;
    reg [7:0] z4209_assgn42090;
    reg [7:0] z1211_assgn1211;
    wire [7:0] c1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4213_assgn4213;
    reg [7:0] z4213_assgn42130;
    reg [7:0] z1213_assgn1213;
    wire [7:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4217_assgn4217;
    reg [7:0] z4217_assgn42170;
    reg [7:0] z1215_assgn1215;
    wire [7:0] d1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4233_assgn4233;
    reg [7:0] z4233_assgn42330;
    reg [7:0] z1229_assgn1229;
    wire [7:0] b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4237_assgn4237;
    reg [7:0] z4237_assgn42370;
    reg [7:0] z1231_assgn1231;
    wire [7:0] b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4243_assgn4243;
    reg [7:0] z4243_assgn42430;
    reg [7:0] z4243_assgn42431;
    reg [7:0] z1235_assgn1235;
    wire [7:0] i1_hpc10_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] axorb_1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4249_assgn4249;
    reg [7:0] z4249_assgn42490;
    reg [7:0] z4249_assgn42491;
    reg [7:0] z1239_assgn1239;
    wire [7:0] i2_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_hpc10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_hpc10_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4265_assgn4265;
    reg [7:0] z4265_assgn42650;
    reg [7:0] z1253_assgn1253;
    wire [7:0] b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4269_assgn4269;
    reg [7:0] z4269_assgn42690;
    reg [7:0] z1255_assgn1255;
    wire [7:0] b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] a0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4275_assgn4275;
    reg [7:0] z4275_assgn42750;
    reg [7:0] z4275_assgn42751;
    reg [7:0] z1259_assgn1259;
    wire [7:0] i1_hpc11_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] a1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4281_assgn4281;
    reg [7:0] z4281_assgn42810;
    reg [7:0] z4281_assgn42811;
    reg [7:0] z1263_assgn1263;
    wire [7:0] i2_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_hpc11_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_hpc11_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4301_assgn4301;
    reg [7:0] z4301_assgn43010;
    reg [7:0] z1281_assgn1281;
    wire [7:0] b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4305_assgn4305;
    reg [7:0] z4305_assgn43050;
    reg [7:0] z1283_assgn1283;
    wire [7:0] b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] b0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4311_assgn4311;
    reg [7:0] z4311_assgn43110;
    reg [7:0] z4311_assgn43111;
    reg [7:0] z1287_assgn1287;
    wire [7:0] i1_hpc12_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] b1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4317_assgn4317;
    reg [7:0] z4317_assgn43170;
    reg [7:0] z4317_assgn43171;
    reg [7:0] z1291_assgn1291;
    wire [7:0] i2_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_hpc12_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_hpc12_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4333_assgn4333;
    reg [7:0] z4333_assgn43330;
    reg [7:0] z4333_assgn43331;
    reg [7:0] z4333_assgn43332;
    reg [7:0] z1305_assgn1305;
    wire [7:0] p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4337_assgn4337;
    reg [7:0] z4337_assgn43370;
    reg [7:0] z4337_assgn43371;
    reg [7:0] z4337_assgn43372;
    reg [7:0] z1307_assgn1307;
    wire [7:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G16_inv0_G256_inv0;
    wire [7:0] d1_G16_inv0_G256_inv0;
    wire [7:0] z4345_assgn4345;
    reg [7:0] z4345_assgn43450;
    reg [7:0] z1314_assgn1314;
    wire [7:0] c0xord0_G16_inv0_G256_inv0;
    wire [7:0] z4349_assgn4349;
    reg [7:0] z4349_assgn43490;
    reg [7:0] z1316_assgn1316;
    wire [7:0] c1xord1_G16_inv0_G256_inv0;
    wire [7:0] z4353_assgn4353;
    reg [7:0] z4353_assgn43530;
    reg [7:0] z4353_assgn43531;
    reg [7:0] z4353_assgn43532;
    reg [7:0] z1317_assgn1317;
    wire [7:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4357_assgn4357;
    reg [7:0] z4357_assgn43570;
    reg [7:0] z4357_assgn43571;
    reg [7:0] z4357_assgn43572;
    reg [7:0] z1319_assgn1319;
    wire [7:0] a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4361_assgn4361;
    reg [7:0] z4361_assgn43610;
    reg [7:0] z4361_assgn43611;
    reg [7:0] z4361_assgn43612;
    reg [7:0] z1321_assgn1321;
    wire [7:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4365_assgn4365;
    reg [7:0] z4365_assgn43650;
    reg [7:0] z4365_assgn43651;
    reg [7:0] z4365_assgn43652;
    reg [7:0] z1323_assgn1323;
    wire [7:0] a1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4369_assgn4369;
    reg [7:0] z4369_assgn43690;
    reg [7:0] z4369_assgn43691;
    reg [7:0] z4369_assgn43692;
    reg [7:0] z1325_assgn1325;
    wire [7:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4373_assgn4373;
    reg [7:0] z4373_assgn43730;
    reg [7:0] z4373_assgn43731;
    reg [7:0] z4373_assgn43732;
    reg [7:0] z1327_assgn1327;
    wire [7:0] b1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4377_assgn4377;
    reg [7:0] z4377_assgn43770;
    reg [7:0] z4377_assgn43771;
    reg [7:0] z4377_assgn43772;
    reg [7:0] z1329_assgn1329;
    wire [7:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4381_assgn4381;
    reg [7:0] z4381_assgn43810;
    reg [7:0] z4381_assgn43811;
    reg [7:0] z4381_assgn43812;
    reg [7:0] z1331_assgn1331;
    wire [7:0] b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] e0_G16_inv0_G256_inv0;
    wire [7:0] e1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4401_assgn4401;
    reg [7:0] z4401_assgn44010;
    reg [7:0] z4401_assgn44011;
    reg [7:0] z4401_assgn44012;
    reg [7:0] z1349_assgn1349;
    wire [7:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4405_assgn4405;
    reg [7:0] z4405_assgn44050;
    reg [7:0] z4405_assgn44051;
    reg [7:0] z4405_assgn44052;
    reg [7:0] z1351_assgn1351;
    wire [7:0] a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4409_assgn4409;
    reg [7:0] z4409_assgn44090;
    reg [7:0] z4409_assgn44091;
    reg [7:0] z4409_assgn44092;
    reg [7:0] z1353_assgn1353;
    wire [7:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4413_assgn4413;
    reg [7:0] z4413_assgn44130;
    reg [7:0] z4413_assgn44131;
    reg [7:0] z4413_assgn44132;
    reg [7:0] z1355_assgn1355;
    wire [7:0] a1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4417_assgn4417;
    reg [7:0] z4417_assgn44170;
    reg [7:0] z4417_assgn44171;
    reg [7:0] z4417_assgn44172;
    reg [7:0] z1357_assgn1357;
    wire [7:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4421_assgn4421;
    reg [7:0] z4421_assgn44210;
    reg [7:0] z4421_assgn44211;
    reg [7:0] z4421_assgn44212;
    reg [7:0] z1359_assgn1359;
    wire [7:0] b1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4425_assgn4425;
    reg [7:0] z4425_assgn44250;
    reg [7:0] z1361_assgn1361;
    wire [7:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4429_assgn4429;
    reg [7:0] z4429_assgn44290;
    reg [7:0] z1363_assgn1363;
    wire [7:0] c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4433_assgn4433;
    reg [7:0] z4433_assgn44330;
    reg [7:0] z1365_assgn1365;
    wire [7:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4437_assgn4437;
    reg [7:0] z4437_assgn44370;
    reg [7:0] z1367_assgn1367;
    wire [7:0] c1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4441_assgn4441;
    reg [7:0] z4441_assgn44410;
    reg [7:0] z1369_assgn1369;
    wire [7:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4445_assgn4445;
    reg [7:0] z4445_assgn44450;
    reg [7:0] z1371_assgn1371;
    wire [7:0] d1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4461_assgn4461;
    reg [7:0] z4461_assgn44610;
    reg [7:0] z1385_assgn1385;
    wire [7:0] b0_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4465_assgn4465;
    reg [7:0] z4465_assgn44650;
    reg [7:0] z1387_assgn1387;
    wire [7:0] b1_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4469_assgn4469;
    reg [7:0] z4469_assgn44690;
    reg [7:0] z1389_assgn1389;
    wire [7:0] p2_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4473_assgn4473;
    reg [7:0] z4473_assgn44730;
    reg [7:0] z4473_assgn44731;
    reg [7:0] z4473_assgn44732;
    reg [7:0] z1391_assgn1391;
    wire [7:0] i1_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4477_assgn4477;
    reg [7:0] z4477_assgn44770;
    reg [7:0] z1393_assgn1393;
    wire [7:0] p3_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4481_assgn4481;
    reg [7:0] z4481_assgn44810;
    reg [7:0] z4481_assgn44811;
    reg [7:0] z4481_assgn44812;
    reg [7:0] z1395_assgn1395;
    wire [7:0] i2_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4485_assgn4485;
    reg [7:0] z4485_assgn44850;
    reg [7:0] z1397_assgn1397;
    wire [7:0] p1_hpc10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4489_assgn4489;
    reg [7:0] z4489_assgn44890;
    reg [7:0] z1399_assgn1399;
    wire [7:0] p4_hpc10_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4501_assgn4501;
    reg [7:0] z4501_assgn45010;
    reg [7:0] z1409_assgn1409;
    wire [7:0] b0_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4505_assgn4505;
    reg [7:0] z4505_assgn45050;
    reg [7:0] z1411_assgn1411;
    wire [7:0] b1_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4509_assgn4509;
    reg [7:0] z4509_assgn45090;
    reg [7:0] z1413_assgn1413;
    wire [7:0] p2_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4513_assgn4513;
    reg [7:0] z4513_assgn45130;
    reg [7:0] z4513_assgn45131;
    reg [7:0] z4513_assgn45132;
    reg [7:0] z1415_assgn1415;
    wire [7:0] i1_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4517_assgn4517;
    reg [7:0] z4517_assgn45170;
    reg [7:0] z1417_assgn1417;
    wire [7:0] p3_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4521_assgn4521;
    reg [7:0] z4521_assgn45210;
    reg [7:0] z4521_assgn45211;
    reg [7:0] z4521_assgn45212;
    reg [7:0] z1419_assgn1419;
    wire [7:0] i2_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4525_assgn4525;
    reg [7:0] z4525_assgn45250;
    reg [7:0] z1421_assgn1421;
    wire [7:0] p1_hpc11_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4529_assgn4529;
    reg [7:0] z4529_assgn45290;
    reg [7:0] z1423_assgn1423;
    wire [7:0] p4_hpc11_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4545_assgn4545;
    reg [7:0] z4545_assgn45450;
    reg [7:0] z1437_assgn1437;
    wire [7:0] b0_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4549_assgn4549;
    reg [7:0] z4549_assgn45490;
    reg [7:0] z1439_assgn1439;
    wire [7:0] b1_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4553_assgn4553;
    reg [7:0] z4553_assgn45530;
    reg [7:0] z1441_assgn1441;
    wire [7:0] p2_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4557_assgn4557;
    reg [7:0] z4557_assgn45570;
    reg [7:0] z4557_assgn45571;
    reg [7:0] z4557_assgn45572;
    reg [7:0] z1443_assgn1443;
    wire [7:0] i1_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4561_assgn4561;
    reg [7:0] z4561_assgn45610;
    reg [7:0] z1445_assgn1445;
    wire [7:0] p3_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4565_assgn4565;
    reg [7:0] z4565_assgn45650;
    reg [7:0] z4565_assgn45651;
    reg [7:0] z4565_assgn45652;
    reg [7:0] z1447_assgn1447;
    wire [7:0] i2_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4569_assgn4569;
    reg [7:0] z4569_assgn45690;
    reg [7:0] z1449_assgn1449;
    wire [7:0] p1_hpc12_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4573_assgn4573;
    reg [7:0] z4573_assgn45730;
    reg [7:0] z1451_assgn1451;
    wire [7:0] p4_hpc12_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4585_assgn4585;
    reg [7:0] z4585_assgn45850;
    reg [7:0] z4585_assgn45851;
    reg [7:0] z4585_assgn45852;
    reg [7:0] z4585_assgn45853;
    reg [7:0] z1461_assgn1461;
    wire [7:0] p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4589_assgn4589;
    reg [7:0] z4589_assgn45890;
    reg [7:0] z4589_assgn45891;
    reg [7:0] z4589_assgn45892;
    reg [7:0] z4589_assgn45893;
    reg [7:0] z1463_assgn1463;
    wire [7:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G16_inv0_G256_inv0;
    wire [7:0] p1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4609_assgn4609;
    reg [7:0] z4609_assgn46090;
    reg [7:0] z4609_assgn46091;
    reg [7:0] z4609_assgn46092;
    reg [7:0] z1481_assgn1481;
    wire [7:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4613_assgn4613;
    reg [7:0] z4613_assgn46130;
    reg [7:0] z4613_assgn46131;
    reg [7:0] z4613_assgn46132;
    reg [7:0] z1483_assgn1483;
    wire [7:0] a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4617_assgn4617;
    reg [7:0] z4617_assgn46170;
    reg [7:0] z4617_assgn46171;
    reg [7:0] z4617_assgn46172;
    reg [7:0] z1485_assgn1485;
    wire [7:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4621_assgn4621;
    reg [7:0] z4621_assgn46210;
    reg [7:0] z4621_assgn46211;
    reg [7:0] z4621_assgn46212;
    reg [7:0] z1487_assgn1487;
    wire [7:0] a1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4625_assgn4625;
    reg [7:0] z4625_assgn46250;
    reg [7:0] z4625_assgn46251;
    reg [7:0] z4625_assgn46252;
    reg [7:0] z1489_assgn1489;
    wire [7:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4629_assgn4629;
    reg [7:0] z4629_assgn46290;
    reg [7:0] z4629_assgn46291;
    reg [7:0] z4629_assgn46292;
    reg [7:0] z1491_assgn1491;
    wire [7:0] b1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4633_assgn4633;
    reg [7:0] z4633_assgn46330;
    reg [7:0] z1493_assgn1493;
    wire [7:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4637_assgn4637;
    reg [7:0] z4637_assgn46370;
    reg [7:0] z1495_assgn1495;
    wire [7:0] c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4641_assgn4641;
    reg [7:0] z4641_assgn46410;
    reg [7:0] z1497_assgn1497;
    wire [7:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4645_assgn4645;
    reg [7:0] z4645_assgn46450;
    reg [7:0] z1499_assgn1499;
    wire [7:0] c1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4649_assgn4649;
    reg [7:0] z4649_assgn46490;
    reg [7:0] z1501_assgn1501;
    wire [7:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4653_assgn4653;
    reg [7:0] z4653_assgn46530;
    reg [7:0] z1503_assgn1503;
    wire [7:0] d1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4669_assgn4669;
    reg [7:0] z4669_assgn46690;
    reg [7:0] z1517_assgn1517;
    wire [7:0] b0_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4673_assgn4673;
    reg [7:0] z4673_assgn46730;
    reg [7:0] z1519_assgn1519;
    wire [7:0] b1_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4677_assgn4677;
    reg [7:0] z4677_assgn46770;
    reg [7:0] z1521_assgn1521;
    wire [7:0] p2_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4681_assgn4681;
    reg [7:0] z4681_assgn46810;
    reg [7:0] z4681_assgn46811;
    reg [7:0] z4681_assgn46812;
    reg [7:0] z1523_assgn1523;
    wire [7:0] i1_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4685_assgn4685;
    reg [7:0] z4685_assgn46850;
    reg [7:0] z1525_assgn1525;
    wire [7:0] p3_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4689_assgn4689;
    reg [7:0] z4689_assgn46890;
    reg [7:0] z4689_assgn46891;
    reg [7:0] z4689_assgn46892;
    reg [7:0] z1527_assgn1527;
    wire [7:0] i2_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4693_assgn4693;
    reg [7:0] z4693_assgn46930;
    reg [7:0] z1529_assgn1529;
    wire [7:0] p1_hpc10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4697_assgn4697;
    reg [7:0] z4697_assgn46970;
    reg [7:0] z1531_assgn1531;
    wire [7:0] p4_hpc10_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4709_assgn4709;
    reg [7:0] z4709_assgn47090;
    reg [7:0] z1541_assgn1541;
    wire [7:0] b0_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4713_assgn4713;
    reg [7:0] z4713_assgn47130;
    reg [7:0] z1543_assgn1543;
    wire [7:0] b1_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4717_assgn4717;
    reg [7:0] z4717_assgn47170;
    reg [7:0] z1545_assgn1545;
    wire [7:0] p2_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4721_assgn4721;
    reg [7:0] z4721_assgn47210;
    reg [7:0] z4721_assgn47211;
    reg [7:0] z4721_assgn47212;
    reg [7:0] z1547_assgn1547;
    wire [7:0] i1_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4725_assgn4725;
    reg [7:0] z4725_assgn47250;
    reg [7:0] z1549_assgn1549;
    wire [7:0] p3_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4729_assgn4729;
    reg [7:0] z4729_assgn47290;
    reg [7:0] z4729_assgn47291;
    reg [7:0] z4729_assgn47292;
    reg [7:0] z1551_assgn1551;
    wire [7:0] i2_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4733_assgn4733;
    reg [7:0] z4733_assgn47330;
    reg [7:0] z1553_assgn1553;
    wire [7:0] p1_hpc11_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4737_assgn4737;
    reg [7:0] z4737_assgn47370;
    reg [7:0] z1555_assgn1555;
    wire [7:0] p4_hpc11_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4753_assgn4753;
    reg [7:0] z4753_assgn47530;
    reg [7:0] z1569_assgn1569;
    wire [7:0] b0_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4757_assgn4757;
    reg [7:0] z4757_assgn47570;
    reg [7:0] z1571_assgn1571;
    wire [7:0] b1_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4761_assgn4761;
    reg [7:0] z4761_assgn47610;
    reg [7:0] z1573_assgn1573;
    wire [7:0] p2_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4765_assgn4765;
    reg [7:0] z4765_assgn47650;
    reg [7:0] z4765_assgn47651;
    reg [7:0] z4765_assgn47652;
    reg [7:0] z1575_assgn1575;
    wire [7:0] i1_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4769_assgn4769;
    reg [7:0] z4769_assgn47690;
    reg [7:0] z1577_assgn1577;
    wire [7:0] p3_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4773_assgn4773;
    reg [7:0] z4773_assgn47730;
    reg [7:0] z4773_assgn47731;
    reg [7:0] z4773_assgn47732;
    reg [7:0] z1579_assgn1579;
    wire [7:0] i2_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4777_assgn4777;
    reg [7:0] z4777_assgn47770;
    reg [7:0] z1581_assgn1581;
    wire [7:0] p1_hpc12_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4781_assgn4781;
    reg [7:0] z4781_assgn47810;
    reg [7:0] z1583_assgn1583;
    wire [7:0] p4_hpc12_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4793_assgn4793;
    reg [7:0] z4793_assgn47930;
    reg [7:0] z4793_assgn47931;
    reg [7:0] z4793_assgn47932;
    reg [7:0] z4793_assgn47933;
    reg [7:0] z1593_assgn1593;
    wire [7:0] p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4797_assgn4797;
    reg [7:0] z4797_assgn47970;
    reg [7:0] z4797_assgn47971;
    reg [7:0] z4797_assgn47972;
    reg [7:0] z4797_assgn47973;
    reg [7:0] z1595_assgn1595;
    wire [7:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G16_inv0_G256_inv0;
    wire [7:0] q1_G16_inv0_G256_inv0;
    wire [7:0] z4805_assgn4805;
    reg [7:0] z4805_assgn48050;
    reg [7:0] z4805_assgn48051;
    reg [7:0] z4805_assgn48052;
    reg [7:0] z4805_assgn48053;
    reg [7:0] z1601_assgn1601;
    wire [7:0] p0ls2_G16_inv0_G256_inv0;
    wire [7:0] z4809_assgn4809;
    reg [7:0] z4809_assgn48090;
    reg [7:0] z4809_assgn48091;
    reg [7:0] z4809_assgn48092;
    reg [7:0] z4809_assgn48093;
    reg [7:0] z1603_assgn1603;
    wire [7:0] p1ls2_G16_inv0_G256_inv0;
    wire [7:0] e0_G256_inv0;
    wire [7:0] e1_G256_inv0;
    wire [7:0] r00_G16_mul1_G256_inv0;
    wire [7:0] v_r1_G16_mul1_G256_inv0;
    wire [7:0] r20_G16_mul1_G256_inv0;
    wire [7:0] r30_G16_mul1_G256_inv0;
    wire [7:0] r40_G16_mul1_G256_inv0;
    wire [7:0] r50_G16_mul1_G256_inv0;
    wire [7:0] r60_G16_mul1_G256_inv0;
    wire [7:0] r70_G16_mul1_G256_inv0;
    wire [7:0] r80_G16_mul1_G256_inv0;
    wire [7:0] r90_G16_mul1_G256_inv0;
    wire [7:0] r100_G16_mul1_G256_inv0;
    wire [7:0] r110_G16_mul1_G256_inv0;
    wire [7:0] r120_G16_mul1_G256_inv0;
    wire [7:0] r130_G16_mul1_G256_inv0;
    wire [7:0] r140_G16_mul1_G256_inv0;
    wire [7:0] r150_G16_mul1_G256_inv0;
    wire [7:0] r160_G16_mul1_G256_inv0;
    wire [7:0] r170_G16_mul1_G256_inv0;
    wire [7:0] z4853_assgn4853;
    reg [7:0] z4853_assgn48530;
    reg [7:0] z4853_assgn48531;
    reg [7:0] z4853_assgn48532;
    reg [7:0] z4853_assgn48533;
    reg [7:0] z1645_assgn1645;
    wire [7:0] a0_0_G16_mul1_G256_inv0;
    wire [7:0] z4857_assgn4857;
    reg [7:0] z4857_assgn48570;
    reg [7:0] z4857_assgn48571;
    reg [7:0] z4857_assgn48572;
    reg [7:0] z4857_assgn48573;
    reg [7:0] z1647_assgn1647;
    wire [7:0] a1_0_G16_mul1_G256_inv0;
    wire [7:0] z4861_assgn4861;
    reg [7:0] z4861_assgn48610;
    reg [7:0] z4861_assgn48611;
    reg [7:0] z4861_assgn48612;
    reg [7:0] z4861_assgn48613;
    reg [7:0] z1649_assgn1649;
    wire [7:0] a0_G16_mul1_G256_inv0;
    wire [7:0] z4865_assgn4865;
    reg [7:0] z4865_assgn48650;
    reg [7:0] z4865_assgn48651;
    reg [7:0] z4865_assgn48652;
    reg [7:0] z4865_assgn48653;
    reg [7:0] z1651_assgn1651;
    wire [7:0] a1_G16_mul1_G256_inv0;
    wire [7:0] z4869_assgn4869;
    reg [7:0] z4869_assgn48690;
    reg [7:0] z4869_assgn48691;
    reg [7:0] z4869_assgn48692;
    reg [7:0] z4869_assgn48693;
    reg [7:0] z1653_assgn1653;
    wire [7:0] b0_G16_mul1_G256_inv0;
    wire [7:0] z4873_assgn4873;
    reg [7:0] z4873_assgn48730;
    reg [7:0] z4873_assgn48731;
    reg [7:0] z4873_assgn48732;
    reg [7:0] z4873_assgn48733;
    reg [7:0] z1655_assgn1655;
    wire [7:0] b1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G16_mul1_G256_inv0;
    wire [7:0] c0_G16_mul1_G256_inv0;
    wire [7:0] c1_G16_mul1_G256_inv0;
    wire [7:0] d0_G16_mul1_G256_inv0;
    wire [7:0] d1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4909_assgn4909;
    reg [7:0] z4909_assgn49090;
    reg [7:0] z4909_assgn49091;
    reg [7:0] z4909_assgn49092;
    reg [7:0] z4909_assgn49093;
    reg [7:0] z1689_assgn1689;
    wire [7:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4913_assgn4913;
    reg [7:0] z4913_assgn49130;
    reg [7:0] z4913_assgn49131;
    reg [7:0] z4913_assgn49132;
    reg [7:0] z4913_assgn49133;
    reg [7:0] z1691_assgn1691;
    wire [7:0] a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4917_assgn4917;
    reg [7:0] z4917_assgn49170;
    reg [7:0] z4917_assgn49171;
    reg [7:0] z4917_assgn49172;
    reg [7:0] z4917_assgn49173;
    reg [7:0] z1693_assgn1693;
    wire [7:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4921_assgn4921;
    reg [7:0] z4921_assgn49210;
    reg [7:0] z4921_assgn49211;
    reg [7:0] z4921_assgn49212;
    reg [7:0] z4921_assgn49213;
    reg [7:0] z1695_assgn1695;
    wire [7:0] a1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4925_assgn4925;
    reg [7:0] z4925_assgn49250;
    reg [7:0] z4925_assgn49251;
    reg [7:0] z4925_assgn49252;
    reg [7:0] z4925_assgn49253;
    reg [7:0] z1697_assgn1697;
    wire [7:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4929_assgn4929;
    reg [7:0] z4929_assgn49290;
    reg [7:0] z4929_assgn49291;
    reg [7:0] z4929_assgn49292;
    reg [7:0] z4929_assgn49293;
    reg [7:0] z1699_assgn1699;
    wire [7:0] b1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4961_assgn4961;
    reg [7:0] z4961_assgn49610;
    reg [7:0] z4961_assgn49611;
    reg [7:0] z4961_assgn49612;
    reg [7:0] z4961_assgn49613;
    reg [7:0] z1729_assgn1729;
    wire [7:0] p2_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4965_assgn4965;
    reg [7:0] z4965_assgn49650;
    reg [7:0] z4965_assgn49651;
    reg [7:0] z4965_assgn49652;
    reg [7:0] z4965_assgn49653;
    reg [7:0] z1731_assgn1731;
    wire [7:0] i1_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4969_assgn4969;
    reg [7:0] z4969_assgn49690;
    reg [7:0] z4969_assgn49691;
    reg [7:0] z4969_assgn49692;
    reg [7:0] z4969_assgn49693;
    reg [7:0] z1733_assgn1733;
    wire [7:0] p3_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4973_assgn4973;
    reg [7:0] z4973_assgn49730;
    reg [7:0] z4973_assgn49731;
    reg [7:0] z4973_assgn49732;
    reg [7:0] z4973_assgn49733;
    reg [7:0] z1735_assgn1735;
    wire [7:0] i2_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4977_assgn4977;
    reg [7:0] z4977_assgn49770;
    reg [7:0] z4977_assgn49771;
    reg [7:0] z4977_assgn49772;
    reg [7:0] z4977_assgn49773;
    reg [7:0] z1737_assgn1737;
    wire [7:0] p1_hpc10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4981_assgn4981;
    reg [7:0] z4981_assgn49810;
    reg [7:0] z4981_assgn49811;
    reg [7:0] z4981_assgn49812;
    reg [7:0] z4981_assgn49813;
    reg [7:0] z1739_assgn1739;
    wire [7:0] p4_hpc10_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4997_assgn4997;
    reg [7:0] z4997_assgn49970;
    reg [7:0] z4997_assgn49971;
    reg [7:0] z4997_assgn49972;
    reg [7:0] z4997_assgn49973;
    reg [7:0] z1753_assgn1753;
    wire [7:0] p2_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5001_assgn5001;
    reg [7:0] z5001_assgn50010;
    reg [7:0] z5001_assgn50011;
    reg [7:0] z5001_assgn50012;
    reg [7:0] z5001_assgn50013;
    reg [7:0] z1755_assgn1755;
    wire [7:0] i1_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5005_assgn5005;
    reg [7:0] z5005_assgn50050;
    reg [7:0] z5005_assgn50051;
    reg [7:0] z5005_assgn50052;
    reg [7:0] z5005_assgn50053;
    reg [7:0] z1757_assgn1757;
    wire [7:0] p3_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5009_assgn5009;
    reg [7:0] z5009_assgn50090;
    reg [7:0] z5009_assgn50091;
    reg [7:0] z5009_assgn50092;
    reg [7:0] z5009_assgn50093;
    reg [7:0] z1759_assgn1759;
    wire [7:0] i2_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5013_assgn5013;
    reg [7:0] z5013_assgn50130;
    reg [7:0] z5013_assgn50131;
    reg [7:0] z5013_assgn50132;
    reg [7:0] z5013_assgn50133;
    reg [7:0] z1761_assgn1761;
    wire [7:0] p1_hpc11_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5017_assgn5017;
    reg [7:0] z5017_assgn50170;
    reg [7:0] z5017_assgn50171;
    reg [7:0] z5017_assgn50172;
    reg [7:0] z5017_assgn50173;
    reg [7:0] z1763_assgn1763;
    wire [7:0] p4_hpc11_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5037_assgn5037;
    reg [7:0] z5037_assgn50370;
    reg [7:0] z5037_assgn50371;
    reg [7:0] z5037_assgn50372;
    reg [7:0] z5037_assgn50373;
    reg [7:0] z1781_assgn1781;
    wire [7:0] p2_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5041_assgn5041;
    reg [7:0] z5041_assgn50410;
    reg [7:0] z5041_assgn50411;
    reg [7:0] z5041_assgn50412;
    reg [7:0] z5041_assgn50413;
    reg [7:0] z1783_assgn1783;
    wire [7:0] i1_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5045_assgn5045;
    reg [7:0] z5045_assgn50450;
    reg [7:0] z5045_assgn50451;
    reg [7:0] z5045_assgn50452;
    reg [7:0] z5045_assgn50453;
    reg [7:0] z1785_assgn1785;
    wire [7:0] p3_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5049_assgn5049;
    reg [7:0] z5049_assgn50490;
    reg [7:0] z5049_assgn50491;
    reg [7:0] z5049_assgn50492;
    reg [7:0] z5049_assgn50493;
    reg [7:0] z1787_assgn1787;
    wire [7:0] i2_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5053_assgn5053;
    reg [7:0] z5053_assgn50530;
    reg [7:0] z5053_assgn50531;
    reg [7:0] z5053_assgn50532;
    reg [7:0] z5053_assgn50533;
    reg [7:0] z1789_assgn1789;
    wire [7:0] p1_hpc12_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5057_assgn5057;
    reg [7:0] z5057_assgn50570;
    reg [7:0] z5057_assgn50571;
    reg [7:0] z5057_assgn50572;
    reg [7:0] z5057_assgn50573;
    reg [7:0] z1791_assgn1791;
    wire [7:0] p4_hpc12_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5069_assgn5069;
    reg [7:0] z5069_assgn50690;
    reg [7:0] z5069_assgn50691;
    reg [7:0] z5069_assgn50692;
    reg [7:0] z5069_assgn50693;
    reg [7:0] z5069_assgn50694;
    reg [7:0] z1801_assgn1801;
    wire [7:0] p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5073_assgn5073;
    reg [7:0] z5073_assgn50730;
    reg [7:0] z5073_assgn50731;
    reg [7:0] z5073_assgn50732;
    reg [7:0] z5073_assgn50733;
    reg [7:0] z5073_assgn50734;
    reg [7:0] z1803_assgn1803;
    wire [7:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G16_mul1_G256_inv0;
    wire [7:0] e1_G16_mul1_G256_inv0;
    wire [7:0] z5081_assgn5081;
    reg [7:0] z5081_assgn50810;
    reg [7:0] z5081_assgn50811;
    reg [7:0] z5081_assgn50812;
    reg [7:0] z5081_assgn50813;
    reg [7:0] z5081_assgn50814;
    reg [7:0] z1809_assgn1809;
    wire [7:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5085_assgn5085;
    reg [7:0] z5085_assgn50850;
    reg [7:0] z5085_assgn50851;
    reg [7:0] z5085_assgn50852;
    reg [7:0] z5085_assgn50853;
    reg [7:0] z5085_assgn50854;
    reg [7:0] z1811_assgn1811;
    wire [7:0] a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5089_assgn5089;
    reg [7:0] z5089_assgn50890;
    reg [7:0] z5089_assgn50891;
    reg [7:0] z5089_assgn50892;
    reg [7:0] z5089_assgn50893;
    reg [7:0] z5089_assgn50894;
    reg [7:0] z1813_assgn1813;
    wire [7:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5093_assgn5093;
    reg [7:0] z5093_assgn50930;
    reg [7:0] z5093_assgn50931;
    reg [7:0] z5093_assgn50932;
    reg [7:0] z5093_assgn50933;
    reg [7:0] z5093_assgn50934;
    reg [7:0] z1815_assgn1815;
    wire [7:0] a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5097_assgn5097;
    reg [7:0] z5097_assgn50970;
    reg [7:0] z5097_assgn50971;
    reg [7:0] z5097_assgn50972;
    reg [7:0] z5097_assgn50973;
    reg [7:0] z5097_assgn50974;
    reg [7:0] z1817_assgn1817;
    wire [7:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5101_assgn5101;
    reg [7:0] z5101_assgn51010;
    reg [7:0] z5101_assgn51011;
    reg [7:0] z5101_assgn51012;
    reg [7:0] z5101_assgn51013;
    reg [7:0] z5101_assgn51014;
    reg [7:0] z1819_assgn1819;
    wire [7:0] b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5113_assgn5113;
    reg [7:0] z5113_assgn51130;
    reg [7:0] z5113_assgn51131;
    reg [7:0] z5113_assgn51132;
    reg [7:0] z5113_assgn51133;
    reg [7:0] z5113_assgn51134;
    reg [7:0] z1829_assgn1829;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5117_assgn5117;
    reg [7:0] z5117_assgn51170;
    reg [7:0] z5117_assgn51171;
    reg [7:0] z5117_assgn51172;
    reg [7:0] z5117_assgn51173;
    reg [7:0] z5117_assgn51174;
    reg [7:0] z1831_assgn1831;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] e01_G16_mul1_G256_inv0;
    wire [7:0] e11_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5137_assgn5137;
    reg [7:0] z5137_assgn51370;
    reg [7:0] z5137_assgn51371;
    reg [7:0] z5137_assgn51372;
    reg [7:0] z5137_assgn51373;
    reg [7:0] z1849_assgn1849;
    wire [7:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5141_assgn5141;
    reg [7:0] z5141_assgn51410;
    reg [7:0] z5141_assgn51411;
    reg [7:0] z5141_assgn51412;
    reg [7:0] z5141_assgn51413;
    reg [7:0] z1851_assgn1851;
    wire [7:0] a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5145_assgn5145;
    reg [7:0] z5145_assgn51450;
    reg [7:0] z5145_assgn51451;
    reg [7:0] z5145_assgn51452;
    reg [7:0] z5145_assgn51453;
    reg [7:0] z1853_assgn1853;
    wire [7:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5149_assgn5149;
    reg [7:0] z5149_assgn51490;
    reg [7:0] z5149_assgn51491;
    reg [7:0] z5149_assgn51492;
    reg [7:0] z5149_assgn51493;
    reg [7:0] z1855_assgn1855;
    wire [7:0] a1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5153_assgn5153;
    reg [7:0] z5153_assgn51530;
    reg [7:0] z5153_assgn51531;
    reg [7:0] z5153_assgn51532;
    reg [7:0] z5153_assgn51533;
    reg [7:0] z1857_assgn1857;
    wire [7:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5157_assgn5157;
    reg [7:0] z5157_assgn51570;
    reg [7:0] z5157_assgn51571;
    reg [7:0] z5157_assgn51572;
    reg [7:0] z5157_assgn51573;
    reg [7:0] z1859_assgn1859;
    wire [7:0] b1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5189_assgn5189;
    reg [7:0] z5189_assgn51890;
    reg [7:0] z5189_assgn51891;
    reg [7:0] z5189_assgn51892;
    reg [7:0] z5189_assgn51893;
    reg [7:0] z1889_assgn1889;
    wire [7:0] p2_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5193_assgn5193;
    reg [7:0] z5193_assgn51930;
    reg [7:0] z5193_assgn51931;
    reg [7:0] z5193_assgn51932;
    reg [7:0] z5193_assgn51933;
    reg [7:0] z1891_assgn1891;
    wire [7:0] i1_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5197_assgn5197;
    reg [7:0] z5197_assgn51970;
    reg [7:0] z5197_assgn51971;
    reg [7:0] z5197_assgn51972;
    reg [7:0] z5197_assgn51973;
    reg [7:0] z1893_assgn1893;
    wire [7:0] p3_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5201_assgn5201;
    reg [7:0] z5201_assgn52010;
    reg [7:0] z5201_assgn52011;
    reg [7:0] z5201_assgn52012;
    reg [7:0] z5201_assgn52013;
    reg [7:0] z1895_assgn1895;
    wire [7:0] i2_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5205_assgn5205;
    reg [7:0] z5205_assgn52050;
    reg [7:0] z5205_assgn52051;
    reg [7:0] z5205_assgn52052;
    reg [7:0] z5205_assgn52053;
    reg [7:0] z1897_assgn1897;
    wire [7:0] p1_hpc10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5209_assgn5209;
    reg [7:0] z5209_assgn52090;
    reg [7:0] z5209_assgn52091;
    reg [7:0] z5209_assgn52092;
    reg [7:0] z5209_assgn52093;
    reg [7:0] z1899_assgn1899;
    wire [7:0] p4_hpc10_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5225_assgn5225;
    reg [7:0] z5225_assgn52250;
    reg [7:0] z5225_assgn52251;
    reg [7:0] z5225_assgn52252;
    reg [7:0] z5225_assgn52253;
    reg [7:0] z1913_assgn1913;
    wire [7:0] p2_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5229_assgn5229;
    reg [7:0] z5229_assgn52290;
    reg [7:0] z5229_assgn52291;
    reg [7:0] z5229_assgn52292;
    reg [7:0] z5229_assgn52293;
    reg [7:0] z1915_assgn1915;
    wire [7:0] i1_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5233_assgn5233;
    reg [7:0] z5233_assgn52330;
    reg [7:0] z5233_assgn52331;
    reg [7:0] z5233_assgn52332;
    reg [7:0] z5233_assgn52333;
    reg [7:0] z1917_assgn1917;
    wire [7:0] p3_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5237_assgn5237;
    reg [7:0] z5237_assgn52370;
    reg [7:0] z5237_assgn52371;
    reg [7:0] z5237_assgn52372;
    reg [7:0] z5237_assgn52373;
    reg [7:0] z1919_assgn1919;
    wire [7:0] i2_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5241_assgn5241;
    reg [7:0] z5241_assgn52410;
    reg [7:0] z5241_assgn52411;
    reg [7:0] z5241_assgn52412;
    reg [7:0] z5241_assgn52413;
    reg [7:0] z1921_assgn1921;
    wire [7:0] p1_hpc11_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5245_assgn5245;
    reg [7:0] z5245_assgn52450;
    reg [7:0] z5245_assgn52451;
    reg [7:0] z5245_assgn52452;
    reg [7:0] z5245_assgn52453;
    reg [7:0] z1923_assgn1923;
    wire [7:0] p4_hpc11_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5265_assgn5265;
    reg [7:0] z5265_assgn52650;
    reg [7:0] z5265_assgn52651;
    reg [7:0] z5265_assgn52652;
    reg [7:0] z5265_assgn52653;
    reg [7:0] z1941_assgn1941;
    wire [7:0] p2_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5269_assgn5269;
    reg [7:0] z5269_assgn52690;
    reg [7:0] z5269_assgn52691;
    reg [7:0] z5269_assgn52692;
    reg [7:0] z5269_assgn52693;
    reg [7:0] z1943_assgn1943;
    wire [7:0] i1_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5273_assgn5273;
    reg [7:0] z5273_assgn52730;
    reg [7:0] z5273_assgn52731;
    reg [7:0] z5273_assgn52732;
    reg [7:0] z5273_assgn52733;
    reg [7:0] z1945_assgn1945;
    wire [7:0] p3_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5277_assgn5277;
    reg [7:0] z5277_assgn52770;
    reg [7:0] z5277_assgn52771;
    reg [7:0] z5277_assgn52772;
    reg [7:0] z5277_assgn52773;
    reg [7:0] z1947_assgn1947;
    wire [7:0] i2_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5281_assgn5281;
    reg [7:0] z5281_assgn52810;
    reg [7:0] z5281_assgn52811;
    reg [7:0] z5281_assgn52812;
    reg [7:0] z5281_assgn52813;
    reg [7:0] z1949_assgn1949;
    wire [7:0] p1_hpc12_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5285_assgn5285;
    reg [7:0] z5285_assgn52850;
    reg [7:0] z5285_assgn52851;
    reg [7:0] z5285_assgn52852;
    reg [7:0] z5285_assgn52853;
    reg [7:0] z1951_assgn1951;
    wire [7:0] p4_hpc12_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5297_assgn5297;
    reg [7:0] z5297_assgn52970;
    reg [7:0] z5297_assgn52971;
    reg [7:0] z5297_assgn52972;
    reg [7:0] z5297_assgn52973;
    reg [7:0] z5297_assgn52974;
    reg [7:0] z1961_assgn1961;
    wire [7:0] p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5301_assgn5301;
    reg [7:0] z5301_assgn53010;
    reg [7:0] z5301_assgn53011;
    reg [7:0] z5301_assgn53012;
    reg [7:0] z5301_assgn53013;
    reg [7:0] z5301_assgn53014;
    reg [7:0] z1963_assgn1963;
    wire [7:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G16_mul1_G256_inv0;
    wire [7:0] p0_G16_mul1_G256_inv0;
    wire [7:0] p1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5325_assgn5325;
    reg [7:0] z5325_assgn53250;
    reg [7:0] z5325_assgn53251;
    reg [7:0] z5325_assgn53252;
    reg [7:0] z5325_assgn53253;
    reg [7:0] z1985_assgn1985;
    wire [7:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5329_assgn5329;
    reg [7:0] z5329_assgn53290;
    reg [7:0] z5329_assgn53291;
    reg [7:0] z5329_assgn53292;
    reg [7:0] z5329_assgn53293;
    reg [7:0] z1987_assgn1987;
    wire [7:0] a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5333_assgn5333;
    reg [7:0] z5333_assgn53330;
    reg [7:0] z5333_assgn53331;
    reg [7:0] z5333_assgn53332;
    reg [7:0] z5333_assgn53333;
    reg [7:0] z1989_assgn1989;
    wire [7:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5337_assgn5337;
    reg [7:0] z5337_assgn53370;
    reg [7:0] z5337_assgn53371;
    reg [7:0] z5337_assgn53372;
    reg [7:0] z5337_assgn53373;
    reg [7:0] z1991_assgn1991;
    wire [7:0] a1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5341_assgn5341;
    reg [7:0] z5341_assgn53410;
    reg [7:0] z5341_assgn53411;
    reg [7:0] z5341_assgn53412;
    reg [7:0] z5341_assgn53413;
    reg [7:0] z1993_assgn1993;
    wire [7:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5345_assgn5345;
    reg [7:0] z5345_assgn53450;
    reg [7:0] z5345_assgn53451;
    reg [7:0] z5345_assgn53452;
    reg [7:0] z5345_assgn53453;
    reg [7:0] z1995_assgn1995;
    wire [7:0] b1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5377_assgn5377;
    reg [7:0] z5377_assgn53770;
    reg [7:0] z5377_assgn53771;
    reg [7:0] z5377_assgn53772;
    reg [7:0] z5377_assgn53773;
    reg [7:0] z2025_assgn2025;
    wire [7:0] p2_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5381_assgn5381;
    reg [7:0] z5381_assgn53810;
    reg [7:0] z5381_assgn53811;
    reg [7:0] z5381_assgn53812;
    reg [7:0] z5381_assgn53813;
    reg [7:0] z2027_assgn2027;
    wire [7:0] i1_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5385_assgn5385;
    reg [7:0] z5385_assgn53850;
    reg [7:0] z5385_assgn53851;
    reg [7:0] z5385_assgn53852;
    reg [7:0] z5385_assgn53853;
    reg [7:0] z2029_assgn2029;
    wire [7:0] p3_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5389_assgn5389;
    reg [7:0] z5389_assgn53890;
    reg [7:0] z5389_assgn53891;
    reg [7:0] z5389_assgn53892;
    reg [7:0] z5389_assgn53893;
    reg [7:0] z2031_assgn2031;
    wire [7:0] i2_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5393_assgn5393;
    reg [7:0] z5393_assgn53930;
    reg [7:0] z5393_assgn53931;
    reg [7:0] z5393_assgn53932;
    reg [7:0] z5393_assgn53933;
    reg [7:0] z2033_assgn2033;
    wire [7:0] p1_hpc10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5397_assgn5397;
    reg [7:0] z5397_assgn53970;
    reg [7:0] z5397_assgn53971;
    reg [7:0] z5397_assgn53972;
    reg [7:0] z5397_assgn53973;
    reg [7:0] z2035_assgn2035;
    wire [7:0] p4_hpc10_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5413_assgn5413;
    reg [7:0] z5413_assgn54130;
    reg [7:0] z5413_assgn54131;
    reg [7:0] z5413_assgn54132;
    reg [7:0] z5413_assgn54133;
    reg [7:0] z2049_assgn2049;
    wire [7:0] p2_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5417_assgn5417;
    reg [7:0] z5417_assgn54170;
    reg [7:0] z5417_assgn54171;
    reg [7:0] z5417_assgn54172;
    reg [7:0] z5417_assgn54173;
    reg [7:0] z2051_assgn2051;
    wire [7:0] i1_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5421_assgn5421;
    reg [7:0] z5421_assgn54210;
    reg [7:0] z5421_assgn54211;
    reg [7:0] z5421_assgn54212;
    reg [7:0] z5421_assgn54213;
    reg [7:0] z2053_assgn2053;
    wire [7:0] p3_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5425_assgn5425;
    reg [7:0] z5425_assgn54250;
    reg [7:0] z5425_assgn54251;
    reg [7:0] z5425_assgn54252;
    reg [7:0] z5425_assgn54253;
    reg [7:0] z2055_assgn2055;
    wire [7:0] i2_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5429_assgn5429;
    reg [7:0] z5429_assgn54290;
    reg [7:0] z5429_assgn54291;
    reg [7:0] z5429_assgn54292;
    reg [7:0] z5429_assgn54293;
    reg [7:0] z2057_assgn2057;
    wire [7:0] p1_hpc11_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5433_assgn5433;
    reg [7:0] z5433_assgn54330;
    reg [7:0] z5433_assgn54331;
    reg [7:0] z5433_assgn54332;
    reg [7:0] z5433_assgn54333;
    reg [7:0] z2059_assgn2059;
    wire [7:0] p4_hpc11_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5453_assgn5453;
    reg [7:0] z5453_assgn54530;
    reg [7:0] z5453_assgn54531;
    reg [7:0] z5453_assgn54532;
    reg [7:0] z5453_assgn54533;
    reg [7:0] z2077_assgn2077;
    wire [7:0] p2_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5457_assgn5457;
    reg [7:0] z5457_assgn54570;
    reg [7:0] z5457_assgn54571;
    reg [7:0] z5457_assgn54572;
    reg [7:0] z5457_assgn54573;
    reg [7:0] z2079_assgn2079;
    wire [7:0] i1_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5461_assgn5461;
    reg [7:0] z5461_assgn54610;
    reg [7:0] z5461_assgn54611;
    reg [7:0] z5461_assgn54612;
    reg [7:0] z5461_assgn54613;
    reg [7:0] z2081_assgn2081;
    wire [7:0] p3_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5465_assgn5465;
    reg [7:0] z5465_assgn54650;
    reg [7:0] z5465_assgn54651;
    reg [7:0] z5465_assgn54652;
    reg [7:0] z5465_assgn54653;
    reg [7:0] z2083_assgn2083;
    wire [7:0] i2_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5469_assgn5469;
    reg [7:0] z5469_assgn54690;
    reg [7:0] z5469_assgn54691;
    reg [7:0] z5469_assgn54692;
    reg [7:0] z5469_assgn54693;
    reg [7:0] z2085_assgn2085;
    wire [7:0] p1_hpc12_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5473_assgn5473;
    reg [7:0] z5473_assgn54730;
    reg [7:0] z5473_assgn54731;
    reg [7:0] z5473_assgn54732;
    reg [7:0] z5473_assgn54733;
    reg [7:0] z2087_assgn2087;
    wire [7:0] p4_hpc12_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5485_assgn5485;
    reg [7:0] z5485_assgn54850;
    reg [7:0] z5485_assgn54851;
    reg [7:0] z5485_assgn54852;
    reg [7:0] z5485_assgn54853;
    reg [7:0] z5485_assgn54854;
    reg [7:0] z2097_assgn2097;
    wire [7:0] p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5489_assgn5489;
    reg [7:0] z5489_assgn54890;
    reg [7:0] z5489_assgn54891;
    reg [7:0] z5489_assgn54892;
    reg [7:0] z5489_assgn54893;
    reg [7:0] z5489_assgn54894;
    reg [7:0] z2099_assgn2099;
    wire [7:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G16_mul1_G256_inv0;
    wire [7:0] q0_G16_mul1_G256_inv0;
    wire [7:0] q1_G16_mul1_G256_inv0;
    wire [7:0] z5501_assgn5501;
    reg [7:0] z5501_assgn55010;
    reg [7:0] z5501_assgn55011;
    reg [7:0] z5501_assgn55012;
    reg [7:0] z5501_assgn55013;
    reg [7:0] z5501_assgn55014;
    reg [7:0] z2109_assgn2109;
    wire [7:0] p0ls2_G16_mul1_G256_inv0;
    wire [7:0] z5505_assgn5505;
    reg [7:0] z5505_assgn55050;
    reg [7:0] z5505_assgn55051;
    reg [7:0] z5505_assgn55052;
    reg [7:0] z5505_assgn55053;
    reg [7:0] z5505_assgn55054;
    reg [7:0] z2111_assgn2111;
    wire [7:0] p1ls2_G16_mul1_G256_inv0;
    wire [7:0] p0_G256_inv0;
    wire [7:0] p1_G256_inv0;
    wire [7:0] r00_G16_mul2_G256_inv0;
    wire [7:0] v_r1_G16_mul2_G256_inv0;
    wire [7:0] r20_G16_mul2_G256_inv0;
    wire [7:0] r30_G16_mul2_G256_inv0;
    wire [7:0] r40_G16_mul2_G256_inv0;
    wire [7:0] r50_G16_mul2_G256_inv0;
    wire [7:0] r60_G16_mul2_G256_inv0;
    wire [7:0] r70_G16_mul2_G256_inv0;
    wire [7:0] r80_G16_mul2_G256_inv0;
    wire [7:0] r90_G16_mul2_G256_inv0;
    wire [7:0] r100_G16_mul2_G256_inv0;
    wire [7:0] r110_G16_mul2_G256_inv0;
    wire [7:0] r120_G16_mul2_G256_inv0;
    wire [7:0] r130_G16_mul2_G256_inv0;
    wire [7:0] r140_G16_mul2_G256_inv0;
    wire [7:0] r150_G16_mul2_G256_inv0;
    wire [7:0] r160_G16_mul2_G256_inv0;
    wire [7:0] r170_G16_mul2_G256_inv0;
    wire [7:0] z5549_assgn5549;
    reg [7:0] z5549_assgn55490;
    reg [7:0] z5549_assgn55491;
    reg [7:0] z5549_assgn55492;
    reg [7:0] z5549_assgn55493;
    reg [7:0] z2153_assgn2153;
    wire [7:0] a0_0_G16_mul2_G256_inv0;
    wire [7:0] z5553_assgn5553;
    reg [7:0] z5553_assgn55530;
    reg [7:0] z5553_assgn55531;
    reg [7:0] z5553_assgn55532;
    reg [7:0] z5553_assgn55533;
    reg [7:0] z2155_assgn2155;
    wire [7:0] a1_0_G16_mul2_G256_inv0;
    wire [7:0] z5557_assgn5557;
    reg [7:0] z5557_assgn55570;
    reg [7:0] z5557_assgn55571;
    reg [7:0] z5557_assgn55572;
    reg [7:0] z5557_assgn55573;
    reg [7:0] z2157_assgn2157;
    wire [7:0] a0_G16_mul2_G256_inv0;
    wire [7:0] z5561_assgn5561;
    reg [7:0] z5561_assgn55610;
    reg [7:0] z5561_assgn55611;
    reg [7:0] z5561_assgn55612;
    reg [7:0] z5561_assgn55613;
    reg [7:0] z2159_assgn2159;
    wire [7:0] a1_G16_mul2_G256_inv0;
    wire [7:0] z5565_assgn5565;
    reg [7:0] z5565_assgn55650;
    reg [7:0] z5565_assgn55651;
    reg [7:0] z5565_assgn55652;
    reg [7:0] z5565_assgn55653;
    reg [7:0] z2161_assgn2161;
    wire [7:0] b0_G16_mul2_G256_inv0;
    wire [7:0] z5569_assgn5569;
    reg [7:0] z5569_assgn55690;
    reg [7:0] z5569_assgn55691;
    reg [7:0] z5569_assgn55692;
    reg [7:0] z5569_assgn55693;
    reg [7:0] z2163_assgn2163;
    wire [7:0] b1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G16_mul2_G256_inv0;
    wire [7:0] c0_G16_mul2_G256_inv0;
    wire [7:0] c1_G16_mul2_G256_inv0;
    wire [7:0] d0_G16_mul2_G256_inv0;
    wire [7:0] d1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5605_assgn5605;
    reg [7:0] z5605_assgn56050;
    reg [7:0] z5605_assgn56051;
    reg [7:0] z5605_assgn56052;
    reg [7:0] z5605_assgn56053;
    reg [7:0] z2197_assgn2197;
    wire [7:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5609_assgn5609;
    reg [7:0] z5609_assgn56090;
    reg [7:0] z5609_assgn56091;
    reg [7:0] z5609_assgn56092;
    reg [7:0] z5609_assgn56093;
    reg [7:0] z2199_assgn2199;
    wire [7:0] a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5613_assgn5613;
    reg [7:0] z5613_assgn56130;
    reg [7:0] z5613_assgn56131;
    reg [7:0] z5613_assgn56132;
    reg [7:0] z5613_assgn56133;
    reg [7:0] z2201_assgn2201;
    wire [7:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5617_assgn5617;
    reg [7:0] z5617_assgn56170;
    reg [7:0] z5617_assgn56171;
    reg [7:0] z5617_assgn56172;
    reg [7:0] z5617_assgn56173;
    reg [7:0] z2203_assgn2203;
    wire [7:0] a1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5621_assgn5621;
    reg [7:0] z5621_assgn56210;
    reg [7:0] z5621_assgn56211;
    reg [7:0] z5621_assgn56212;
    reg [7:0] z5621_assgn56213;
    reg [7:0] z2205_assgn2205;
    wire [7:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5625_assgn5625;
    reg [7:0] z5625_assgn56250;
    reg [7:0] z5625_assgn56251;
    reg [7:0] z5625_assgn56252;
    reg [7:0] z5625_assgn56253;
    reg [7:0] z2207_assgn2207;
    wire [7:0] b1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5657_assgn5657;
    reg [7:0] z5657_assgn56570;
    reg [7:0] z5657_assgn56571;
    reg [7:0] z5657_assgn56572;
    reg [7:0] z5657_assgn56573;
    reg [7:0] z2237_assgn2237;
    wire [7:0] p2_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5661_assgn5661;
    reg [7:0] z5661_assgn56610;
    reg [7:0] z5661_assgn56611;
    reg [7:0] z5661_assgn56612;
    reg [7:0] z5661_assgn56613;
    reg [7:0] z2239_assgn2239;
    wire [7:0] i1_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5665_assgn5665;
    reg [7:0] z5665_assgn56650;
    reg [7:0] z5665_assgn56651;
    reg [7:0] z5665_assgn56652;
    reg [7:0] z5665_assgn56653;
    reg [7:0] z2241_assgn2241;
    wire [7:0] p3_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5669_assgn5669;
    reg [7:0] z5669_assgn56690;
    reg [7:0] z5669_assgn56691;
    reg [7:0] z5669_assgn56692;
    reg [7:0] z5669_assgn56693;
    reg [7:0] z2243_assgn2243;
    wire [7:0] i2_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5673_assgn5673;
    reg [7:0] z5673_assgn56730;
    reg [7:0] z5673_assgn56731;
    reg [7:0] z5673_assgn56732;
    reg [7:0] z5673_assgn56733;
    reg [7:0] z2245_assgn2245;
    wire [7:0] p1_hpc10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5677_assgn5677;
    reg [7:0] z5677_assgn56770;
    reg [7:0] z5677_assgn56771;
    reg [7:0] z5677_assgn56772;
    reg [7:0] z5677_assgn56773;
    reg [7:0] z2247_assgn2247;
    wire [7:0] p4_hpc10_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5693_assgn5693;
    reg [7:0] z5693_assgn56930;
    reg [7:0] z5693_assgn56931;
    reg [7:0] z5693_assgn56932;
    reg [7:0] z5693_assgn56933;
    reg [7:0] z2261_assgn2261;
    wire [7:0] p2_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5697_assgn5697;
    reg [7:0] z5697_assgn56970;
    reg [7:0] z5697_assgn56971;
    reg [7:0] z5697_assgn56972;
    reg [7:0] z5697_assgn56973;
    reg [7:0] z2263_assgn2263;
    wire [7:0] i1_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5701_assgn5701;
    reg [7:0] z5701_assgn57010;
    reg [7:0] z5701_assgn57011;
    reg [7:0] z5701_assgn57012;
    reg [7:0] z5701_assgn57013;
    reg [7:0] z2265_assgn2265;
    wire [7:0] p3_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5705_assgn5705;
    reg [7:0] z5705_assgn57050;
    reg [7:0] z5705_assgn57051;
    reg [7:0] z5705_assgn57052;
    reg [7:0] z5705_assgn57053;
    reg [7:0] z2267_assgn2267;
    wire [7:0] i2_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5709_assgn5709;
    reg [7:0] z5709_assgn57090;
    reg [7:0] z5709_assgn57091;
    reg [7:0] z5709_assgn57092;
    reg [7:0] z5709_assgn57093;
    reg [7:0] z2269_assgn2269;
    wire [7:0] p1_hpc11_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5713_assgn5713;
    reg [7:0] z5713_assgn57130;
    reg [7:0] z5713_assgn57131;
    reg [7:0] z5713_assgn57132;
    reg [7:0] z5713_assgn57133;
    reg [7:0] z2271_assgn2271;
    wire [7:0] p4_hpc11_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5733_assgn5733;
    reg [7:0] z5733_assgn57330;
    reg [7:0] z5733_assgn57331;
    reg [7:0] z5733_assgn57332;
    reg [7:0] z5733_assgn57333;
    reg [7:0] z2289_assgn2289;
    wire [7:0] p2_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5737_assgn5737;
    reg [7:0] z5737_assgn57370;
    reg [7:0] z5737_assgn57371;
    reg [7:0] z5737_assgn57372;
    reg [7:0] z5737_assgn57373;
    reg [7:0] z2291_assgn2291;
    wire [7:0] i1_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5741_assgn5741;
    reg [7:0] z5741_assgn57410;
    reg [7:0] z5741_assgn57411;
    reg [7:0] z5741_assgn57412;
    reg [7:0] z5741_assgn57413;
    reg [7:0] z2293_assgn2293;
    wire [7:0] p3_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5745_assgn5745;
    reg [7:0] z5745_assgn57450;
    reg [7:0] z5745_assgn57451;
    reg [7:0] z5745_assgn57452;
    reg [7:0] z5745_assgn57453;
    reg [7:0] z2295_assgn2295;
    wire [7:0] i2_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5749_assgn5749;
    reg [7:0] z5749_assgn57490;
    reg [7:0] z5749_assgn57491;
    reg [7:0] z5749_assgn57492;
    reg [7:0] z5749_assgn57493;
    reg [7:0] z2297_assgn2297;
    wire [7:0] p1_hpc12_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5753_assgn5753;
    reg [7:0] z5753_assgn57530;
    reg [7:0] z5753_assgn57531;
    reg [7:0] z5753_assgn57532;
    reg [7:0] z5753_assgn57533;
    reg [7:0] z2299_assgn2299;
    wire [7:0] p4_hpc12_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5765_assgn5765;
    reg [7:0] z5765_assgn57650;
    reg [7:0] z5765_assgn57651;
    reg [7:0] z5765_assgn57652;
    reg [7:0] z5765_assgn57653;
    reg [7:0] z5765_assgn57654;
    reg [7:0] z2309_assgn2309;
    wire [7:0] p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5769_assgn5769;
    reg [7:0] z5769_assgn57690;
    reg [7:0] z5769_assgn57691;
    reg [7:0] z5769_assgn57692;
    reg [7:0] z5769_assgn57693;
    reg [7:0] z5769_assgn57694;
    reg [7:0] z2311_assgn2311;
    wire [7:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G16_mul2_G256_inv0;
    wire [7:0] e1_G16_mul2_G256_inv0;
    wire [7:0] z5777_assgn5777;
    reg [7:0] z5777_assgn57770;
    reg [7:0] z5777_assgn57771;
    reg [7:0] z5777_assgn57772;
    reg [7:0] z5777_assgn57773;
    reg [7:0] z5777_assgn57774;
    reg [7:0] z2317_assgn2317;
    wire [7:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5781_assgn5781;
    reg [7:0] z5781_assgn57810;
    reg [7:0] z5781_assgn57811;
    reg [7:0] z5781_assgn57812;
    reg [7:0] z5781_assgn57813;
    reg [7:0] z5781_assgn57814;
    reg [7:0] z2319_assgn2319;
    wire [7:0] a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5785_assgn5785;
    reg [7:0] z5785_assgn57850;
    reg [7:0] z5785_assgn57851;
    reg [7:0] z5785_assgn57852;
    reg [7:0] z5785_assgn57853;
    reg [7:0] z5785_assgn57854;
    reg [7:0] z2321_assgn2321;
    wire [7:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5789_assgn5789;
    reg [7:0] z5789_assgn57890;
    reg [7:0] z5789_assgn57891;
    reg [7:0] z5789_assgn57892;
    reg [7:0] z5789_assgn57893;
    reg [7:0] z5789_assgn57894;
    reg [7:0] z2323_assgn2323;
    wire [7:0] a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5793_assgn5793;
    reg [7:0] z5793_assgn57930;
    reg [7:0] z5793_assgn57931;
    reg [7:0] z5793_assgn57932;
    reg [7:0] z5793_assgn57933;
    reg [7:0] z5793_assgn57934;
    reg [7:0] z2325_assgn2325;
    wire [7:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5797_assgn5797;
    reg [7:0] z5797_assgn57970;
    reg [7:0] z5797_assgn57971;
    reg [7:0] z5797_assgn57972;
    reg [7:0] z5797_assgn57973;
    reg [7:0] z5797_assgn57974;
    reg [7:0] z2327_assgn2327;
    wire [7:0] b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5809_assgn5809;
    reg [7:0] z5809_assgn58090;
    reg [7:0] z5809_assgn58091;
    reg [7:0] z5809_assgn58092;
    reg [7:0] z5809_assgn58093;
    reg [7:0] z5809_assgn58094;
    reg [7:0] z2337_assgn2337;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5813_assgn5813;
    reg [7:0] z5813_assgn58130;
    reg [7:0] z5813_assgn58131;
    reg [7:0] z5813_assgn58132;
    reg [7:0] z5813_assgn58133;
    reg [7:0] z5813_assgn58134;
    reg [7:0] z2339_assgn2339;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] e01_G16_mul2_G256_inv0;
    wire [7:0] e11_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5833_assgn5833;
    reg [7:0] z5833_assgn58330;
    reg [7:0] z5833_assgn58331;
    reg [7:0] z5833_assgn58332;
    reg [7:0] z5833_assgn58333;
    reg [7:0] z2357_assgn2357;
    wire [7:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5837_assgn5837;
    reg [7:0] z5837_assgn58370;
    reg [7:0] z5837_assgn58371;
    reg [7:0] z5837_assgn58372;
    reg [7:0] z5837_assgn58373;
    reg [7:0] z2359_assgn2359;
    wire [7:0] a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5841_assgn5841;
    reg [7:0] z5841_assgn58410;
    reg [7:0] z5841_assgn58411;
    reg [7:0] z5841_assgn58412;
    reg [7:0] z5841_assgn58413;
    reg [7:0] z2361_assgn2361;
    wire [7:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5845_assgn5845;
    reg [7:0] z5845_assgn58450;
    reg [7:0] z5845_assgn58451;
    reg [7:0] z5845_assgn58452;
    reg [7:0] z5845_assgn58453;
    reg [7:0] z2363_assgn2363;
    wire [7:0] a1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5849_assgn5849;
    reg [7:0] z5849_assgn58490;
    reg [7:0] z5849_assgn58491;
    reg [7:0] z5849_assgn58492;
    reg [7:0] z5849_assgn58493;
    reg [7:0] z2365_assgn2365;
    wire [7:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5853_assgn5853;
    reg [7:0] z5853_assgn58530;
    reg [7:0] z5853_assgn58531;
    reg [7:0] z5853_assgn58532;
    reg [7:0] z5853_assgn58533;
    reg [7:0] z2367_assgn2367;
    wire [7:0] b1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5885_assgn5885;
    reg [7:0] z5885_assgn58850;
    reg [7:0] z5885_assgn58851;
    reg [7:0] z5885_assgn58852;
    reg [7:0] z5885_assgn58853;
    reg [7:0] z2397_assgn2397;
    wire [7:0] p2_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5889_assgn5889;
    reg [7:0] z5889_assgn58890;
    reg [7:0] z5889_assgn58891;
    reg [7:0] z5889_assgn58892;
    reg [7:0] z5889_assgn58893;
    reg [7:0] z2399_assgn2399;
    wire [7:0] i1_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5893_assgn5893;
    reg [7:0] z5893_assgn58930;
    reg [7:0] z5893_assgn58931;
    reg [7:0] z5893_assgn58932;
    reg [7:0] z5893_assgn58933;
    reg [7:0] z2401_assgn2401;
    wire [7:0] p3_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5897_assgn5897;
    reg [7:0] z5897_assgn58970;
    reg [7:0] z5897_assgn58971;
    reg [7:0] z5897_assgn58972;
    reg [7:0] z5897_assgn58973;
    reg [7:0] z2403_assgn2403;
    wire [7:0] i2_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5901_assgn5901;
    reg [7:0] z5901_assgn59010;
    reg [7:0] z5901_assgn59011;
    reg [7:0] z5901_assgn59012;
    reg [7:0] z5901_assgn59013;
    reg [7:0] z2405_assgn2405;
    wire [7:0] p1_hpc10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5905_assgn5905;
    reg [7:0] z5905_assgn59050;
    reg [7:0] z5905_assgn59051;
    reg [7:0] z5905_assgn59052;
    reg [7:0] z5905_assgn59053;
    reg [7:0] z2407_assgn2407;
    wire [7:0] p4_hpc10_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5921_assgn5921;
    reg [7:0] z5921_assgn59210;
    reg [7:0] z5921_assgn59211;
    reg [7:0] z5921_assgn59212;
    reg [7:0] z5921_assgn59213;
    reg [7:0] z2421_assgn2421;
    wire [7:0] p2_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5925_assgn5925;
    reg [7:0] z5925_assgn59250;
    reg [7:0] z5925_assgn59251;
    reg [7:0] z5925_assgn59252;
    reg [7:0] z5925_assgn59253;
    reg [7:0] z2423_assgn2423;
    wire [7:0] i1_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5929_assgn5929;
    reg [7:0] z5929_assgn59290;
    reg [7:0] z5929_assgn59291;
    reg [7:0] z5929_assgn59292;
    reg [7:0] z5929_assgn59293;
    reg [7:0] z2425_assgn2425;
    wire [7:0] p3_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5933_assgn5933;
    reg [7:0] z5933_assgn59330;
    reg [7:0] z5933_assgn59331;
    reg [7:0] z5933_assgn59332;
    reg [7:0] z5933_assgn59333;
    reg [7:0] z2427_assgn2427;
    wire [7:0] i2_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5937_assgn5937;
    reg [7:0] z5937_assgn59370;
    reg [7:0] z5937_assgn59371;
    reg [7:0] z5937_assgn59372;
    reg [7:0] z5937_assgn59373;
    reg [7:0] z2429_assgn2429;
    wire [7:0] p1_hpc11_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5941_assgn5941;
    reg [7:0] z5941_assgn59410;
    reg [7:0] z5941_assgn59411;
    reg [7:0] z5941_assgn59412;
    reg [7:0] z5941_assgn59413;
    reg [7:0] z2431_assgn2431;
    wire [7:0] p4_hpc11_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5961_assgn5961;
    reg [7:0] z5961_assgn59610;
    reg [7:0] z5961_assgn59611;
    reg [7:0] z5961_assgn59612;
    reg [7:0] z5961_assgn59613;
    reg [7:0] z2449_assgn2449;
    wire [7:0] p2_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5965_assgn5965;
    reg [7:0] z5965_assgn59650;
    reg [7:0] z5965_assgn59651;
    reg [7:0] z5965_assgn59652;
    reg [7:0] z5965_assgn59653;
    reg [7:0] z2451_assgn2451;
    wire [7:0] i1_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5969_assgn5969;
    reg [7:0] z5969_assgn59690;
    reg [7:0] z5969_assgn59691;
    reg [7:0] z5969_assgn59692;
    reg [7:0] z5969_assgn59693;
    reg [7:0] z2453_assgn2453;
    wire [7:0] p3_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5973_assgn5973;
    reg [7:0] z5973_assgn59730;
    reg [7:0] z5973_assgn59731;
    reg [7:0] z5973_assgn59732;
    reg [7:0] z5973_assgn59733;
    reg [7:0] z2455_assgn2455;
    wire [7:0] i2_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5977_assgn5977;
    reg [7:0] z5977_assgn59770;
    reg [7:0] z5977_assgn59771;
    reg [7:0] z5977_assgn59772;
    reg [7:0] z5977_assgn59773;
    reg [7:0] z2457_assgn2457;
    wire [7:0] p1_hpc12_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5981_assgn5981;
    reg [7:0] z5981_assgn59810;
    reg [7:0] z5981_assgn59811;
    reg [7:0] z5981_assgn59812;
    reg [7:0] z5981_assgn59813;
    reg [7:0] z2459_assgn2459;
    wire [7:0] p4_hpc12_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5993_assgn5993;
    reg [7:0] z5993_assgn59930;
    reg [7:0] z5993_assgn59931;
    reg [7:0] z5993_assgn59932;
    reg [7:0] z5993_assgn59933;
    reg [7:0] z5993_assgn59934;
    reg [7:0] z2469_assgn2469;
    wire [7:0] p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5997_assgn5997;
    reg [7:0] z5997_assgn59970;
    reg [7:0] z5997_assgn59971;
    reg [7:0] z5997_assgn59972;
    reg [7:0] z5997_assgn59973;
    reg [7:0] z5997_assgn59974;
    reg [7:0] z2471_assgn2471;
    wire [7:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G16_mul2_G256_inv0;
    wire [7:0] p0_G16_mul2_G256_inv0;
    wire [7:0] p1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6021_assgn6021;
    reg [7:0] z6021_assgn60210;
    reg [7:0] z6021_assgn60211;
    reg [7:0] z6021_assgn60212;
    reg [7:0] z6021_assgn60213;
    reg [7:0] z2493_assgn2493;
    wire [7:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6025_assgn6025;
    reg [7:0] z6025_assgn60250;
    reg [7:0] z6025_assgn60251;
    reg [7:0] z6025_assgn60252;
    reg [7:0] z6025_assgn60253;
    reg [7:0] z2495_assgn2495;
    wire [7:0] a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6029_assgn6029;
    reg [7:0] z6029_assgn60290;
    reg [7:0] z6029_assgn60291;
    reg [7:0] z6029_assgn60292;
    reg [7:0] z6029_assgn60293;
    reg [7:0] z2497_assgn2497;
    wire [7:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6033_assgn6033;
    reg [7:0] z6033_assgn60330;
    reg [7:0] z6033_assgn60331;
    reg [7:0] z6033_assgn60332;
    reg [7:0] z6033_assgn60333;
    reg [7:0] z2499_assgn2499;
    wire [7:0] a1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6037_assgn6037;
    reg [7:0] z6037_assgn60370;
    reg [7:0] z6037_assgn60371;
    reg [7:0] z6037_assgn60372;
    reg [7:0] z6037_assgn60373;
    reg [7:0] z2501_assgn2501;
    wire [7:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6041_assgn6041;
    reg [7:0] z6041_assgn60410;
    reg [7:0] z6041_assgn60411;
    reg [7:0] z6041_assgn60412;
    reg [7:0] z6041_assgn60413;
    reg [7:0] z2503_assgn2503;
    wire [7:0] b1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6073_assgn6073;
    reg [7:0] z6073_assgn60730;
    reg [7:0] z6073_assgn60731;
    reg [7:0] z6073_assgn60732;
    reg [7:0] z6073_assgn60733;
    reg [7:0] z2533_assgn2533;
    wire [7:0] p2_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6077_assgn6077;
    reg [7:0] z6077_assgn60770;
    reg [7:0] z6077_assgn60771;
    reg [7:0] z6077_assgn60772;
    reg [7:0] z6077_assgn60773;
    reg [7:0] z2535_assgn2535;
    wire [7:0] i1_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6081_assgn6081;
    reg [7:0] z6081_assgn60810;
    reg [7:0] z6081_assgn60811;
    reg [7:0] z6081_assgn60812;
    reg [7:0] z6081_assgn60813;
    reg [7:0] z2537_assgn2537;
    wire [7:0] p3_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6085_assgn6085;
    reg [7:0] z6085_assgn60850;
    reg [7:0] z6085_assgn60851;
    reg [7:0] z6085_assgn60852;
    reg [7:0] z6085_assgn60853;
    reg [7:0] z2539_assgn2539;
    wire [7:0] i2_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6089_assgn6089;
    reg [7:0] z6089_assgn60890;
    reg [7:0] z6089_assgn60891;
    reg [7:0] z6089_assgn60892;
    reg [7:0] z6089_assgn60893;
    reg [7:0] z2541_assgn2541;
    wire [7:0] p1_hpc10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6093_assgn6093;
    reg [7:0] z6093_assgn60930;
    reg [7:0] z6093_assgn60931;
    reg [7:0] z6093_assgn60932;
    reg [7:0] z6093_assgn60933;
    reg [7:0] z2543_assgn2543;
    wire [7:0] p4_hpc10_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc10_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc10_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6109_assgn6109;
    reg [7:0] z6109_assgn61090;
    reg [7:0] z6109_assgn61091;
    reg [7:0] z6109_assgn61092;
    reg [7:0] z6109_assgn61093;
    reg [7:0] z2557_assgn2557;
    wire [7:0] p2_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6113_assgn6113;
    reg [7:0] z6113_assgn61130;
    reg [7:0] z6113_assgn61131;
    reg [7:0] z6113_assgn61132;
    reg [7:0] z6113_assgn61133;
    reg [7:0] z2559_assgn2559;
    wire [7:0] i1_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6117_assgn6117;
    reg [7:0] z6117_assgn61170;
    reg [7:0] z6117_assgn61171;
    reg [7:0] z6117_assgn61172;
    reg [7:0] z6117_assgn61173;
    reg [7:0] z2561_assgn2561;
    wire [7:0] p3_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6121_assgn6121;
    reg [7:0] z6121_assgn61210;
    reg [7:0] z6121_assgn61211;
    reg [7:0] z6121_assgn61212;
    reg [7:0] z6121_assgn61213;
    reg [7:0] z2563_assgn2563;
    wire [7:0] i2_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6125_assgn6125;
    reg [7:0] z6125_assgn61250;
    reg [7:0] z6125_assgn61251;
    reg [7:0] z6125_assgn61252;
    reg [7:0] z6125_assgn61253;
    reg [7:0] z2565_assgn2565;
    wire [7:0] p1_hpc11_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6129_assgn6129;
    reg [7:0] z6129_assgn61290;
    reg [7:0] z6129_assgn61291;
    reg [7:0] z6129_assgn61292;
    reg [7:0] z6129_assgn61293;
    reg [7:0] z2567_assgn2567;
    wire [7:0] p4_hpc11_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc11_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc11_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b0_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b1_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6149_assgn6149;
    reg [7:0] z6149_assgn61490;
    reg [7:0] z6149_assgn61491;
    reg [7:0] z6149_assgn61492;
    reg [7:0] z6149_assgn61493;
    reg [7:0] z2585_assgn2585;
    wire [7:0] p2_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6153_assgn6153;
    reg [7:0] z6153_assgn61530;
    reg [7:0] z6153_assgn61531;
    reg [7:0] z6153_assgn61532;
    reg [7:0] z6153_assgn61533;
    reg [7:0] z2587_assgn2587;
    wire [7:0] i1_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6157_assgn6157;
    reg [7:0] z6157_assgn61570;
    reg [7:0] z6157_assgn61571;
    reg [7:0] z6157_assgn61572;
    reg [7:0] z6157_assgn61573;
    reg [7:0] z2589_assgn2589;
    wire [7:0] p3_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6161_assgn6161;
    reg [7:0] z6161_assgn61610;
    reg [7:0] z6161_assgn61611;
    reg [7:0] z6161_assgn61612;
    reg [7:0] z6161_assgn61613;
    reg [7:0] z2591_assgn2591;
    wire [7:0] i2_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6165_assgn6165;
    reg [7:0] z6165_assgn61650;
    reg [7:0] z6165_assgn61651;
    reg [7:0] z6165_assgn61652;
    reg [7:0] z6165_assgn61653;
    reg [7:0] z2593_assgn2593;
    wire [7:0] p1_hpc12_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6169_assgn6169;
    reg [7:0] z6169_assgn61690;
    reg [7:0] z6169_assgn61691;
    reg [7:0] z6169_assgn61692;
    reg [7:0] z6169_assgn61693;
    reg [7:0] z2595_assgn2595;
    wire [7:0] p4_hpc12_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_hpc12_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_hpc12_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6181_assgn6181;
    reg [7:0] z6181_assgn61810;
    reg [7:0] z6181_assgn61811;
    reg [7:0] z6181_assgn61812;
    reg [7:0] z6181_assgn61813;
    reg [7:0] z6181_assgn61814;
    reg [7:0] z2605_assgn2605;
    wire [7:0] p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6185_assgn6185;
    reg [7:0] z6185_assgn61850;
    reg [7:0] z6185_assgn61851;
    reg [7:0] z6185_assgn61852;
    reg [7:0] z6185_assgn61853;
    reg [7:0] z6185_assgn61854;
    reg [7:0] z2607_assgn2607;
    wire [7:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G16_mul2_G256_inv0;
    wire [7:0] q0_G16_mul2_G256_inv0;
    wire [7:0] q1_G16_mul2_G256_inv0;
    wire [7:0] z6197_assgn6197;
    reg [7:0] z6197_assgn61970;
    reg [7:0] z6197_assgn61971;
    reg [7:0] z6197_assgn61972;
    reg [7:0] z6197_assgn61973;
    reg [7:0] z6197_assgn61974;
    reg [7:0] z2617_assgn2617;
    wire [7:0] p0ls2_G16_mul2_G256_inv0;
    wire [7:0] z6201_assgn6201;
    reg [7:0] z6201_assgn62010;
    reg [7:0] z6201_assgn62011;
    reg [7:0] z6201_assgn62012;
    reg [7:0] z6201_assgn62013;
    reg [7:0] z6201_assgn62014;
    reg [7:0] z2619_assgn2619;
    wire [7:0] p1ls2_G16_mul2_G256_inv0;
    wire [7:0] q0_G256_inv0;
    wire [7:0] q1_G256_inv0;
    wire [7:0] z6209_assgn6209;
    reg [7:0] z6209_assgn62090;
    reg [7:0] z6209_assgn62091;
    reg [7:0] z6209_assgn62092;
    reg [7:0] z6209_assgn62093;
    reg [7:0] z6209_assgn62094;
    reg [7:0] z2625_assgn2625;
    wire [7:0] p0ls4_G256_inv0;
    wire [7:0] z6213_assgn6213;
    reg [7:0] z6213_assgn62130;
    reg [7:0] z6213_assgn62131;
    reg [7:0] z6213_assgn62132;
    reg [7:0] z6213_assgn62133;
    reg [7:0] z6213_assgn62134;
    reg [7:0] z2627_assgn2627;
    wire [7:0] p1ls4_G256_inv0;
    wire [7:0] t4;
    wire [7:0] t5;
    wire [7:0] y_G256_newbasis1;
    wire [7:0] tempy1_G256_newbasis1;
    wire [7:0] z6225_assgn6225;
    reg [7:0] z6225_assgn62250;
    reg [7:0] z6225_assgn62251;
    reg [7:0] z6225_assgn62252;
    reg [7:0] z6225_assgn62253;
    reg [7:0] z6225_assgn62254;
    reg [7:0] z2637_assgn2637;
    wire [7:0] cond1_G256_newbasis1;
    wire [7:0] negCond1_G256_newbasis1;
    wire [7:0] yxorb1_G256_newbasis1;
    wire [7:0] z6233_assgn6233;
    reg [7:0] z6233_assgn62330;
    reg [7:0] z6233_assgn62331;
    reg [7:0] z6233_assgn62332;
    reg [7:0] z6233_assgn62333;
    reg [7:0] z6233_assgn62334;
    reg [7:0] z2643_assgn2643;
    wire [7:0] ny1_G256_newbasis1;
    wire [7:0] z6237_assgn6237;
    reg [7:0] z6237_assgn62370;
    reg [7:0] z6237_assgn62371;
    reg [7:0] z6237_assgn62372;
    reg [7:0] z6237_assgn62373;
    reg [7:0] z6237_assgn62374;
    reg [7:0] z2646_assgn2646;
    wire [7:0] tempyIntoNegCond1_G256_newbasis1;
    wire [7:0] y1_G256_newbasis1;
    wire [7:0] z6243_assgn6243;
    reg [7:0] z6243_assgn62430;
    reg [7:0] z6243_assgn62431;
    reg [7:0] z6243_assgn62432;
    reg [7:0] z6243_assgn62433;
    reg [7:0] z6243_assgn62434;
    reg [7:0] z2649_assgn2649;
    wire [7:0] x1_G256_newbasis1;
    wire [7:0] tempy2_G256_newbasis1;
    wire [7:0] z6249_assgn6249;
    reg [7:0] z6249_assgn62490;
    reg [7:0] z6249_assgn62491;
    reg [7:0] z6249_assgn62492;
    reg [7:0] z6249_assgn62493;
    reg [7:0] z6249_assgn62494;
    reg [7:0] z2653_assgn2653;
    wire [7:0] cond2_G256_newbasis1;
    wire [7:0] negCond2_G256_newbasis1;
    wire [7:0] z6255_assgn6255;
    reg [7:0] z6255_assgn62550;
    reg [7:0] z6255_assgn62551;
    reg [7:0] z6255_assgn62552;
    reg [7:0] z6255_assgn62553;
    reg [7:0] z6255_assgn62554;
    reg [7:0] z2657_assgn2657;
    wire [7:0] yxorb2_G256_newbasis1;
    wire [7:0] ny2_G256_newbasis1;
    wire [7:0] tempyIntoNegCond2_G256_newbasis1;
    wire [7:0] y2_G256_newbasis1;
    wire [7:0] z6265_assgn6265;
    reg [7:0] z6265_assgn62650;
    reg [7:0] z6265_assgn62651;
    reg [7:0] z6265_assgn62652;
    reg [7:0] z6265_assgn62653;
    reg [7:0] z6265_assgn62654;
    reg [7:0] z2665_assgn2665;
    wire [7:0] x2_G256_newbasis1;
    wire [7:0] tempy3_G256_newbasis1;
    wire [7:0] z6271_assgn6271;
    reg [7:0] z6271_assgn62710;
    reg [7:0] z6271_assgn62711;
    reg [7:0] z6271_assgn62712;
    reg [7:0] z6271_assgn62713;
    reg [7:0] z6271_assgn62714;
    reg [7:0] z2669_assgn2669;
    wire [7:0] cond3_G256_newbasis1;
    wire [7:0] negCond3_G256_newbasis1;
    wire [7:0] z6277_assgn6277;
    reg [7:0] z6277_assgn62770;
    reg [7:0] z6277_assgn62771;
    reg [7:0] z6277_assgn62772;
    reg [7:0] z6277_assgn62773;
    reg [7:0] z6277_assgn62774;
    reg [7:0] z2673_assgn2673;
    wire [7:0] yxorb3_G256_newbasis1;
    wire [7:0] ny3_G256_newbasis1;
    wire [7:0] tempyIntoNegCond3_G256_newbasis1;
    wire [7:0] y3_G256_newbasis1;
    wire [7:0] z6287_assgn6287;
    reg [7:0] z6287_assgn62870;
    reg [7:0] z6287_assgn62871;
    reg [7:0] z6287_assgn62872;
    reg [7:0] z6287_assgn62873;
    reg [7:0] z6287_assgn62874;
    reg [7:0] z2681_assgn2681;
    wire [7:0] x3_G256_newbasis1;
    wire [7:0] tempy4_G256_newbasis1;
    wire [7:0] z6293_assgn6293;
    reg [7:0] z6293_assgn62930;
    reg [7:0] z6293_assgn62931;
    reg [7:0] z6293_assgn62932;
    reg [7:0] z6293_assgn62933;
    reg [7:0] z6293_assgn62934;
    reg [7:0] z2685_assgn2685;
    wire [7:0] cond4_G256_newbasis1;
    wire [7:0] negCond4_G256_newbasis1;
    wire [7:0] z6299_assgn6299;
    reg [7:0] z6299_assgn62990;
    reg [7:0] z6299_assgn62991;
    reg [7:0] z6299_assgn62992;
    reg [7:0] z6299_assgn62993;
    reg [7:0] z6299_assgn62994;
    reg [7:0] z2689_assgn2689;
    wire [7:0] yxorb4_G256_newbasis1;
    wire [7:0] ny4_G256_newbasis1;
    wire [7:0] tempyIntoNegCond4_G256_newbasis1;
    wire [7:0] y4_G256_newbasis1;
    wire [7:0] z6309_assgn6309;
    reg [7:0] z6309_assgn63090;
    reg [7:0] z6309_assgn63091;
    reg [7:0] z6309_assgn63092;
    reg [7:0] z6309_assgn63093;
    reg [7:0] z6309_assgn63094;
    reg [7:0] z2697_assgn2697;
    wire [7:0] x4_G256_newbasis1;
    wire [7:0] tempy5_G256_newbasis1;
    wire [7:0] z6315_assgn6315;
    reg [7:0] z6315_assgn63150;
    reg [7:0] z6315_assgn63151;
    reg [7:0] z6315_assgn63152;
    reg [7:0] z6315_assgn63153;
    reg [7:0] z6315_assgn63154;
    reg [7:0] z2701_assgn2701;
    wire [7:0] cond5_G256_newbasis1;
    wire [7:0] negCond5_G256_newbasis1;
    wire [7:0] z6321_assgn6321;
    reg [7:0] z6321_assgn63210;
    reg [7:0] z6321_assgn63211;
    reg [7:0] z6321_assgn63212;
    reg [7:0] z6321_assgn63213;
    reg [7:0] z6321_assgn63214;
    reg [7:0] z2705_assgn2705;
    wire [7:0] yxorb5_G256_newbasis1;
    wire [7:0] ny5_G256_newbasis1;
    wire [7:0] tempyIntoNegCond5_G256_newbasis1;
    wire [7:0] y5_G256_newbasis1;
    wire [7:0] z6331_assgn6331;
    reg [7:0] z6331_assgn63310;
    reg [7:0] z6331_assgn63311;
    reg [7:0] z6331_assgn63312;
    reg [7:0] z6331_assgn63313;
    reg [7:0] z6331_assgn63314;
    reg [7:0] z2713_assgn2713;
    wire [7:0] x5_G256_newbasis1;
    wire [7:0] tempy6_G256_newbasis1;
    wire [7:0] z6337_assgn6337;
    reg [7:0] z6337_assgn63370;
    reg [7:0] z6337_assgn63371;
    reg [7:0] z6337_assgn63372;
    reg [7:0] z6337_assgn63373;
    reg [7:0] z6337_assgn63374;
    reg [7:0] z2717_assgn2717;
    wire [7:0] cond6_G256_newbasis1;
    wire [7:0] negCond6_G256_newbasis1;
    wire [7:0] z6343_assgn6343;
    reg [7:0] z6343_assgn63430;
    reg [7:0] z6343_assgn63431;
    reg [7:0] z6343_assgn63432;
    reg [7:0] z6343_assgn63433;
    reg [7:0] z6343_assgn63434;
    reg [7:0] z2721_assgn2721;
    wire [7:0] yxorb6_G256_newbasis1;
    wire [7:0] ny6_G256_newbasis1;
    wire [7:0] tempyIntoNegCond6_G256_newbasis1;
    wire [7:0] y6_G256_newbasis1;
    wire [7:0] z6353_assgn6353;
    reg [7:0] z6353_assgn63530;
    reg [7:0] z6353_assgn63531;
    reg [7:0] z6353_assgn63532;
    reg [7:0] z6353_assgn63533;
    reg [7:0] z6353_assgn63534;
    reg [7:0] z2729_assgn2729;
    wire [7:0] x6_G256_newbasis1;
    wire [7:0] tempy7_G256_newbasis1;
    wire [7:0] z6359_assgn6359;
    reg [7:0] z6359_assgn63590;
    reg [7:0] z6359_assgn63591;
    reg [7:0] z6359_assgn63592;
    reg [7:0] z6359_assgn63593;
    reg [7:0] z6359_assgn63594;
    reg [7:0] z2733_assgn2733;
    wire [7:0] cond7_G256_newbasis1;
    wire [7:0] negCond7_G256_newbasis1;
    wire [7:0] z6365_assgn6365;
    reg [7:0] z6365_assgn63650;
    reg [7:0] z6365_assgn63651;
    reg [7:0] z6365_assgn63652;
    reg [7:0] z6365_assgn63653;
    reg [7:0] z6365_assgn63654;
    reg [7:0] z2737_assgn2737;
    wire [7:0] yxorb7_G256_newbasis1;
    wire [7:0] ny7_G256_newbasis1;
    wire [7:0] tempyIntoNegCond7_G256_newbasis1;
    wire [7:0] y7_G256_newbasis1;
    wire [7:0] z6375_assgn6375;
    reg [7:0] z6375_assgn63750;
    reg [7:0] z6375_assgn63751;
    reg [7:0] z6375_assgn63752;
    reg [7:0] z6375_assgn63753;
    reg [7:0] z6375_assgn63754;
    reg [7:0] z2745_assgn2745;
    wire [7:0] x7_G256_newbasis1;
    wire [7:0] tempy8_G256_newbasis1;
    wire [7:0] z6381_assgn6381;
    reg [7:0] z6381_assgn63810;
    reg [7:0] z6381_assgn63811;
    reg [7:0] z6381_assgn63812;
    reg [7:0] z6381_assgn63813;
    reg [7:0] z6381_assgn63814;
    reg [7:0] z2749_assgn2749;
    wire [7:0] cond8_G256_newbasis1;
    wire [7:0] negCond8_G256_newbasis1;
    wire [7:0] z6387_assgn6387;
    reg [7:0] z6387_assgn63870;
    reg [7:0] z6387_assgn63871;
    reg [7:0] z6387_assgn63872;
    reg [7:0] z6387_assgn63873;
    reg [7:0] z6387_assgn63874;
    reg [7:0] z2753_assgn2753;
    wire [7:0] yxorb8_G256_newbasis1;
    wire [7:0] ny8_G256_newbasis1;
    wire [7:0] tempyIntoNegCond8_G256_newbasis1;
    wire [7:0] y8_G256_newbasis1;
    wire [7:0] z6397_assgn6397;
    reg [7:0] z6397_assgn63970;
    reg [7:0] z6397_assgn63971;
    reg [7:0] z6397_assgn63972;
    reg [7:0] z6397_assgn63973;
    reg [7:0] z6397_assgn63974;
    reg [7:0] z2761_assgn2761;
    wire [7:0] x8_G256_newbasis1;
    wire [7:0] t6;
    wire [7:0] z_y_G256_newbasis1;
    wire [7:0] z_tempy1_G256_newbasis1;
    wire [7:0] z6407_assgn6407;
    reg [7:0] z6407_assgn64070;
    reg [7:0] z6407_assgn64071;
    reg [7:0] z6407_assgn64072;
    reg [7:0] z6407_assgn64073;
    reg [7:0] z6407_assgn64074;
    reg [7:0] z2769_assgn2769;
    wire [7:0] z_cond1_G256_newbasis1;
    wire [7:0] z_negCond1_G256_newbasis1;
    wire [7:0] z_yxorb1_G256_newbasis1;
    wire [7:0] z6415_assgn6415;
    reg [7:0] z6415_assgn64150;
    reg [7:0] z6415_assgn64151;
    reg [7:0] z6415_assgn64152;
    reg [7:0] z6415_assgn64153;
    reg [7:0] z6415_assgn64154;
    reg [7:0] z2775_assgn2775;
    wire [7:0] z_ny1_G256_newbasis1;
    wire [7:0] z6419_assgn6419;
    reg [7:0] z6419_assgn64190;
    reg [7:0] z6419_assgn64191;
    reg [7:0] z6419_assgn64192;
    reg [7:0] z6419_assgn64193;
    reg [7:0] z6419_assgn64194;
    reg [7:0] z2778_assgn2778;
    wire [7:0] z_tempyIntoNegCond1_G256_newbasis1;
    wire [7:0] z_y1_G256_newbasis1;
    wire [7:0] z6425_assgn6425;
    reg [7:0] z6425_assgn64250;
    reg [7:0] z6425_assgn64251;
    reg [7:0] z6425_assgn64252;
    reg [7:0] z6425_assgn64253;
    reg [7:0] z6425_assgn64254;
    reg [7:0] z2781_assgn2781;
    wire [7:0] z_x1_G256_newbasis1;
    wire [7:0] z_tempy2_G256_newbasis1;
    wire [7:0] z6431_assgn6431;
    reg [7:0] z6431_assgn64310;
    reg [7:0] z6431_assgn64311;
    reg [7:0] z6431_assgn64312;
    reg [7:0] z6431_assgn64313;
    reg [7:0] z6431_assgn64314;
    reg [7:0] z2785_assgn2785;
    wire [7:0] z_cond2_G256_newbasis1;
    wire [7:0] z_negCond2_G256_newbasis1;
    wire [7:0] z6437_assgn6437;
    reg [7:0] z6437_assgn64370;
    reg [7:0] z6437_assgn64371;
    reg [7:0] z6437_assgn64372;
    reg [7:0] z6437_assgn64373;
    reg [7:0] z6437_assgn64374;
    reg [7:0] z2789_assgn2789;
    wire [7:0] z_yxorb2_G256_newbasis1;
    wire [7:0] z_ny2_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond2_G256_newbasis1;
    wire [7:0] z_y2_G256_newbasis1;
    wire [7:0] z6447_assgn6447;
    reg [7:0] z6447_assgn64470;
    reg [7:0] z6447_assgn64471;
    reg [7:0] z6447_assgn64472;
    reg [7:0] z6447_assgn64473;
    reg [7:0] z6447_assgn64474;
    reg [7:0] z2797_assgn2797;
    wire [7:0] z_x2_G256_newbasis1;
    wire [7:0] z_tempy3_G256_newbasis1;
    wire [7:0] z6453_assgn6453;
    reg [7:0] z6453_assgn64530;
    reg [7:0] z6453_assgn64531;
    reg [7:0] z6453_assgn64532;
    reg [7:0] z6453_assgn64533;
    reg [7:0] z6453_assgn64534;
    reg [7:0] z2801_assgn2801;
    wire [7:0] z_cond3_G256_newbasis1;
    wire [7:0] z_negCond3_G256_newbasis1;
    wire [7:0] z6459_assgn6459;
    reg [7:0] z6459_assgn64590;
    reg [7:0] z6459_assgn64591;
    reg [7:0] z6459_assgn64592;
    reg [7:0] z6459_assgn64593;
    reg [7:0] z6459_assgn64594;
    reg [7:0] z2805_assgn2805;
    wire [7:0] z_yxorb3_G256_newbasis1;
    wire [7:0] z_ny3_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond3_G256_newbasis1;
    wire [7:0] z_y3_G256_newbasis1;
    wire [7:0] z6469_assgn6469;
    reg [7:0] z6469_assgn64690;
    reg [7:0] z6469_assgn64691;
    reg [7:0] z6469_assgn64692;
    reg [7:0] z6469_assgn64693;
    reg [7:0] z6469_assgn64694;
    reg [7:0] z2813_assgn2813;
    wire [7:0] z_x3_G256_newbasis1;
    wire [7:0] z_tempy4_G256_newbasis1;
    wire [7:0] z6475_assgn6475;
    reg [7:0] z6475_assgn64750;
    reg [7:0] z6475_assgn64751;
    reg [7:0] z6475_assgn64752;
    reg [7:0] z6475_assgn64753;
    reg [7:0] z6475_assgn64754;
    reg [7:0] z2817_assgn2817;
    wire [7:0] z_cond4_G256_newbasis1;
    wire [7:0] z_negCond4_G256_newbasis1;
    wire [7:0] z6481_assgn6481;
    reg [7:0] z6481_assgn64810;
    reg [7:0] z6481_assgn64811;
    reg [7:0] z6481_assgn64812;
    reg [7:0] z6481_assgn64813;
    reg [7:0] z6481_assgn64814;
    reg [7:0] z2821_assgn2821;
    wire [7:0] z_yxorb4_G256_newbasis1;
    wire [7:0] z_ny4_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond4_G256_newbasis1;
    wire [7:0] z_y4_G256_newbasis1;
    wire [7:0] z6491_assgn6491;
    reg [7:0] z6491_assgn64910;
    reg [7:0] z6491_assgn64911;
    reg [7:0] z6491_assgn64912;
    reg [7:0] z6491_assgn64913;
    reg [7:0] z6491_assgn64914;
    reg [7:0] z2829_assgn2829;
    wire [7:0] z_x4_G256_newbasis1;
    wire [7:0] z_tempy5_G256_newbasis1;
    wire [7:0] z6497_assgn6497;
    reg [7:0] z6497_assgn64970;
    reg [7:0] z6497_assgn64971;
    reg [7:0] z6497_assgn64972;
    reg [7:0] z6497_assgn64973;
    reg [7:0] z6497_assgn64974;
    reg [7:0] z2833_assgn2833;
    wire [7:0] z_cond5_G256_newbasis1;
    wire [7:0] z_negCond5_G256_newbasis1;
    wire [7:0] z6503_assgn6503;
    reg [7:0] z6503_assgn65030;
    reg [7:0] z6503_assgn65031;
    reg [7:0] z6503_assgn65032;
    reg [7:0] z6503_assgn65033;
    reg [7:0] z6503_assgn65034;
    reg [7:0] z2837_assgn2837;
    wire [7:0] z_yxorb5_G256_newbasis1;
    wire [7:0] z_ny5_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond5_G256_newbasis1;
    wire [7:0] z_y5_G256_newbasis1;
    wire [7:0] z6513_assgn6513;
    reg [7:0] z6513_assgn65130;
    reg [7:0] z6513_assgn65131;
    reg [7:0] z6513_assgn65132;
    reg [7:0] z6513_assgn65133;
    reg [7:0] z6513_assgn65134;
    reg [7:0] z2845_assgn2845;
    wire [7:0] z_x5_G256_newbasis1;
    wire [7:0] z_tempy6_G256_newbasis1;
    wire [7:0] z6519_assgn6519;
    reg [7:0] z6519_assgn65190;
    reg [7:0] z6519_assgn65191;
    reg [7:0] z6519_assgn65192;
    reg [7:0] z6519_assgn65193;
    reg [7:0] z6519_assgn65194;
    reg [7:0] z2849_assgn2849;
    wire [7:0] z_cond6_G256_newbasis1;
    wire [7:0] z_negCond6_G256_newbasis1;
    wire [7:0] z6525_assgn6525;
    reg [7:0] z6525_assgn65250;
    reg [7:0] z6525_assgn65251;
    reg [7:0] z6525_assgn65252;
    reg [7:0] z6525_assgn65253;
    reg [7:0] z6525_assgn65254;
    reg [7:0] z2853_assgn2853;
    wire [7:0] z_yxorb6_G256_newbasis1;
    wire [7:0] z_ny6_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond6_G256_newbasis1;
    wire [7:0] z_y6_G256_newbasis1;
    wire [7:0] z6535_assgn6535;
    reg [7:0] z6535_assgn65350;
    reg [7:0] z6535_assgn65351;
    reg [7:0] z6535_assgn65352;
    reg [7:0] z6535_assgn65353;
    reg [7:0] z6535_assgn65354;
    reg [7:0] z2861_assgn2861;
    wire [7:0] z_x6_G256_newbasis1;
    wire [7:0] z_tempy7_G256_newbasis1;
    wire [7:0] z6541_assgn6541;
    reg [7:0] z6541_assgn65410;
    reg [7:0] z6541_assgn65411;
    reg [7:0] z6541_assgn65412;
    reg [7:0] z6541_assgn65413;
    reg [7:0] z6541_assgn65414;
    reg [7:0] z2865_assgn2865;
    wire [7:0] z_cond7_G256_newbasis1;
    wire [7:0] z_negCond7_G256_newbasis1;
    wire [7:0] z6547_assgn6547;
    reg [7:0] z6547_assgn65470;
    reg [7:0] z6547_assgn65471;
    reg [7:0] z6547_assgn65472;
    reg [7:0] z6547_assgn65473;
    reg [7:0] z6547_assgn65474;
    reg [7:0] z2869_assgn2869;
    wire [7:0] z_yxorb7_G256_newbasis1;
    wire [7:0] z_ny7_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond7_G256_newbasis1;
    wire [7:0] z_y7_G256_newbasis1;
    wire [7:0] z6557_assgn6557;
    reg [7:0] z6557_assgn65570;
    reg [7:0] z6557_assgn65571;
    reg [7:0] z6557_assgn65572;
    reg [7:0] z6557_assgn65573;
    reg [7:0] z6557_assgn65574;
    reg [7:0] z2877_assgn2877;
    wire [7:0] z_x7_G256_newbasis1;
    wire [7:0] z_tempy8_G256_newbasis1;
    wire [7:0] z6563_assgn6563;
    reg [7:0] z6563_assgn65630;
    reg [7:0] z6563_assgn65631;
    reg [7:0] z6563_assgn65632;
    reg [7:0] z6563_assgn65633;
    reg [7:0] z6563_assgn65634;
    reg [7:0] z2881_assgn2881;
    wire [7:0] z_cond8_G256_newbasis1;
    wire [7:0] z_negCond8_G256_newbasis1;
    wire [7:0] z6569_assgn6569;
    reg [7:0] z6569_assgn65690;
    reg [7:0] z6569_assgn65691;
    reg [7:0] z6569_assgn65692;
    reg [7:0] z6569_assgn65693;
    reg [7:0] z6569_assgn65694;
    reg [7:0] z2885_assgn2885;
    wire [7:0] z_yxorb8_G256_newbasis1;
    wire [7:0] z_ny8_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond8_G256_newbasis1;
    wire [7:0] z_y8_G256_newbasis1;
    wire [7:0] z6579_assgn6579;
    reg [7:0] z6579_assgn65790;
    reg [7:0] z6579_assgn65791;
    reg [7:0] z6579_assgn65792;
    reg [7:0] z6579_assgn65793;
    reg [7:0] z6579_assgn65794;
    reg [7:0] z2893_assgn2893;
    wire [7:0] z_x8_G256_newbasis1;
    wire [7:0] t7;
    wire [7:0] z6585_assgn6585;
    reg [7:0] z6585_assgn65850;
    reg [7:0] z6585_assgn65851;
    reg [7:0] z6585_assgn65852;
    reg [7:0] z6585_assgn65853;
    reg [7:0] z6585_assgn65854;
    reg [7:0] z2897_assgn2897;


    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign r6_inp = r6;
    assign r7_inp = r7;
    assign r8_inp = r8;
    assign r9_inp = r9;
    assign r10_inp = r10;
    assign r11_inp = r11;
    assign r12_inp = r12;
    assign r13_inp = r13;
    assign r14_inp = r14;
    assign r15_inp = r15;
    assign r16_inp = r16;
    assign r17_inp = r17;
    assign r18_inp = r18;
    assign r19_inp = r19;
    assign r20_inp = r20;
    assign r21_inp = r21;
    assign r22_inp = r22;
    assign r23_inp = r23;
    assign r24_inp = r24;
    assign r25_inp = r25;
    assign r26_inp = r26;
    assign r27_inp = r27;
    assign r28_inp = r28;
    assign r29_inp = r29;
    assign r30_inp = r30;
    assign r31_inp = r31;
    assign r32_inp = r32;
    assign r33_inp = r33;
    assign r34_inp = r34;
    assign r35_inp = r35;
    assign r36_inp = r36;
    assign r37_inp = r37;
    assign r38_inp = r38;
    assign r39_inp = r39;
    assign r40_inp = r40;
    assign r41_inp = r41;
    assign r42_inp = r42;
    assign r43_inp = r43;
    assign r44_inp = r44;
    assign r45_inp = r45;
    assign r46_inp = r46;
    assign r47_inp = r47;
    assign r48_inp = r48;
    assign r49_inp = r49;
    assign r50_inp = r50;
    assign r51_inp = r51;
    assign r52_inp = r52;
    assign r53_inp = r53;
    assign r54_inp = r54;
    assign r55_inp = r55;
    assign r56_inp = r56;
    assign r57_inp = r57;
    assign r58_inp = r58;
    assign r59_inp = r59;
    assign r60_inp = r60;
    assign r61_inp = r61;
    assign r62_inp = r62;
    assign r63_inp = r63;
    assign r64_inp = r64;
    assign r65_inp = r65;
    assign r66_inp = r66;
    assign r67_inp = r67;
    assign r68_inp = r68;
    assign r69_inp = r69;
    assign r70_inp = r70;
    assign r71_inp = r71;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempyIntoNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempyIntoNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempyIntoNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempyIntoNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempyIntoNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempyIntoNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempyIntoNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempyIntoNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0);
    assign z3225_assgn3225 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempyIntoNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempyIntoNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempyIntoNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempyIntoNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempyIntoNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempyIntoNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempyIntoNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempyIntoNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempyIntoNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempyIntoNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempyIntoNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempyIntoNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempyIntoNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempyIntoNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempyIntoNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempyIntoNegCond8_G256_newbasis0);
    assign z3357_assgn3357 = (z_x7_G256_newbasis0 >> dec_1_inp);
    assign t3 = z_y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a1_0_G256_inv0 = (t3 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a1xorb1_G256_inv0 = (a1_G256_inv0 ^ b1_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (r0_inp % dec_16_inp);
    assign v_r1_G16_mul0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul0_G256_inv0 = (r5_inp % dec_16_inp);
    assign r60_G16_mul0_G256_inv0 = (r6_inp % dec_16_inp);
    assign r70_G16_mul0_G256_inv0 = (r7_inp % dec_16_inp);
    assign r80_G16_mul0_G256_inv0 = (r8_inp % dec_16_inp);
    assign r90_G16_mul0_G256_inv0 = (r9_inp % dec_16_inp);
    assign r100_G16_mul0_G256_inv0 = (r10_inp % dec_16_inp);
    assign r110_G16_mul0_G256_inv0 = (r11_inp % dec_16_inp);
    assign r120_G16_mul0_G256_inv0 = (r12_inp % dec_16_inp);
    assign r130_G16_mul0_G256_inv0 = (r13_inp % dec_16_inp);
    assign r140_G16_mul0_G256_inv0 = (r14_inp % dec_16_inp);
    assign r150_G16_mul0_G256_inv0 = (r15_inp % dec_16_inp);
    assign r160_G16_mul0_G256_inv0 = (r16_inp % dec_16_inp);
    assign r170_G16_mul0_G256_inv0 = (r17_inp % dec_16_inp);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (v_r1_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ d1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_hpc10_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul0_G256_inv0);
    assign b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc10_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_hpc10_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc10_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc10_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_hpc10_G4_mul0_G16_mul0_G256_inv0 = (p3_hpc10_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc10_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_hpc10_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (i1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (i2_hpc10_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_hpc10_G4_mul0_G16_mul0_G256_inv0_reg);
    assign r00_hpc11_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul0_G256_inv0);
    assign b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc11_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_hpc11_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc11_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc11_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_hpc11_G4_mul0_G16_mul0_G256_inv0 = (p3_hpc11_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc11_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_hpc11_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (i1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (i2_hpc11_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_hpc11_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_hpc12_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0 = (d0_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul0_G256_inv0);
    assign b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0 = (d1_G4_mul0_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc12_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_hpc12_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc12_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc12_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_hpc12_G4_mul0_G16_mul0_G256_inv0 = (p3_hpc12_G4_mul0_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc12_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_hpc12_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (i1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (i2_hpc12_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_hpc12_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign z3661_assgn3661 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << z761_assgn761);
    assign z3665_assgn3665 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << z763_assgn763);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign z3673_assgn3673 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z769_assgn769);
    assign z3677_assgn3677 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z771_assgn771);
    assign z3681_assgn3681 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> z773_assgn773);
    assign z3685_assgn3685 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> z775_assgn775);
    assign z3689_assgn3689 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z777_assgn777);
    assign z3693_assgn3693 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z779_assgn779);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign z3705_assgn3705 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << z789_assgn789);
    assign z3709_assgn3709 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << z791_assgn791);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r60_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r70_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r80_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul0_G256_inv0 = (r90_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul0_G256_inv0 = (r100_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul0_G256_inv0 = (r110_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ d1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_hpc10_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0 = (cxord_0_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul0_G256_inv0);
    assign b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0 = (cxord_1_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc10_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_hpc10_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc10_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc10_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_hpc10_G4_mul1_G16_mul0_G256_inv0 = (p3_hpc10_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc10_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_hpc10_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (i1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (i2_hpc10_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_hpc10_G4_mul1_G16_mul0_G256_inv0_reg);
    assign r00_hpc11_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul0_G256_inv0);
    assign b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc11_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_hpc11_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc11_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc11_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_hpc11_G4_mul1_G16_mul0_G256_inv0 = (p3_hpc11_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc11_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_hpc11_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (i1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (i2_hpc11_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_hpc11_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_hpc12_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0 = (d0_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul0_G256_inv0);
    assign b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0 = (d1_G4_mul1_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc12_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_hpc12_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc12_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc12_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_hpc12_G4_mul1_G16_mul0_G256_inv0 = (p3_hpc12_G4_mul1_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc12_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_hpc12_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (i1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (i2_hpc12_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_hpc12_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign z3841_assgn3841 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << z921_assgn921);
    assign z3845_assgn3845 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << z923_assgn923);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r120_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r130_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r140_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul0_G256_inv0 = (r150_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul0_G256_inv0 = (r160_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul0_G256_inv0 = (r170_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ d1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_hpc10_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0 = (cxord_0_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul0_G256_inv0);
    assign b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0 = (cxord_1_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc10_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_hpc10_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc10_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc10_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_hpc10_G4_mul2_G16_mul0_G256_inv0 = (p3_hpc10_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc10_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_hpc10_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (i1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (i2_hpc10_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_hpc10_G4_mul2_G16_mul0_G256_inv0_reg);
    assign r00_hpc11_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul0_G256_inv0);
    assign b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc11_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_hpc11_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc11_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc11_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_hpc11_G4_mul2_G16_mul0_G256_inv0 = (p3_hpc11_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc11_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_hpc11_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (i1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (i2_hpc11_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_hpc11_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_hpc12_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0 = (d0_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul0_G256_inv0);
    assign b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0 = (d1_G4_mul2_G16_mul0_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc12_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_hpc12_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc12_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc12_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_hpc12_G4_mul2_G16_mul0_G256_inv0 = (p3_hpc12_G4_mul2_G16_mul0_G256_inv0 ^ r10_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc12_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0_reg & b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_hpc12_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0_reg & b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (i1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (i2_hpc12_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_hpc12_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign z3981_assgn3981 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << z1057_assgn1057);
    assign z3985_assgn3985 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << z1059_assgn1059);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign z3997_assgn3997 = dec_2_inp;
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << z1069_assgn1069);
    assign z4001_assgn4001 = dec_2_inp;
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << z1071_assgn1071);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign z4009_assgn4009 = c0_G256_inv0;
    assign c0xord0_G256_inv0 = (z1078_assgn1078 ^ d0_G256_inv0);
    assign z4013_assgn4013 = c1_G256_inv0;
    assign c1xord1_G256_inv0 = (z1080_assgn1080 ^ d1_G256_inv0);
    assign r00_G16_inv0_G256_inv0 = (r18_inp % dec_16_inp);
    assign v_r1_G16_inv0_G256_inv0 = (r19_inp % dec_16_inp);
    assign r20_G16_inv0_G256_inv0 = (r20_inp % dec_16_inp);
    assign r30_G16_inv0_G256_inv0 = (r21_inp % dec_16_inp);
    assign r40_G16_inv0_G256_inv0 = (r22_inp % dec_16_inp);
    assign r50_G16_inv0_G256_inv0 = (r23_inp % dec_16_inp);
    assign r60_G16_inv0_G256_inv0 = (r24_inp % dec_16_inp);
    assign r70_G16_inv0_G256_inv0 = (r25_inp % dec_16_inp);
    assign r80_G16_inv0_G256_inv0 = (r26_inp % dec_16_inp);
    assign r90_G16_inv0_G256_inv0 = (r27_inp % dec_16_inp);
    assign r100_G16_inv0_G256_inv0 = (r28_inp % dec_16_inp);
    assign r110_G16_inv0_G256_inv0 = (r29_inp % dec_16_inp);
    assign r120_G16_inv0_G256_inv0 = (r30_inp % dec_16_inp);
    assign r130_G16_inv0_G256_inv0 = (r31_inp % dec_16_inp);
    assign r140_G16_inv0_G256_inv0 = (r32_inp % dec_16_inp);
    assign r150_G16_inv0_G256_inv0 = (r33_inp % dec_16_inp);
    assign r160_G16_inv0_G256_inv0 = (r34_inp % dec_16_inp);
    assign r170_G16_inv0_G256_inv0 = (r35_inp % dec_16_inp);
    assign z4053_assgn4053 = dec_12_inp;
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & z1117_assgn1117);
    assign z4057_assgn4057 = dec_12_inp;
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1119_assgn1119);
    assign z4061_assgn4061 = dec_2_inp;
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> z1121_assgn1121);
    assign z4065_assgn4065 = dec_2_inp;
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> z1123_assgn1123);
    assign z4069_assgn4069 = dec_3_inp;
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & z1125_assgn1125);
    assign z4073_assgn4073 = dec_3_inp;
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1127_assgn1127);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a1xorb1_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 ^ b1_G16_inv0_G256_inv0);
    assign z4081_assgn4081 = dec_2_inp;
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1133_assgn1133);
    assign z4085_assgn4085 = dec_2_inp;
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1135_assgn1135);
    assign z4089_assgn4089 = dec_1_inp;
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> z1137_assgn1137);
    assign z4093_assgn4093 = dec_1_inp;
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> z1139_assgn1139);
    assign z4097_assgn4097 = dec_1_inp;
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1141_assgn1141);
    assign z4101_assgn4101 = dec_1_inp;
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1143_assgn1143);
    assign z4105_assgn4105 = dec_1_inp;
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << z1145_assgn1145);
    assign z4109_assgn4109 = dec_1_inp;
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << z1147_assgn1147);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign z4117_assgn4117 = dec_2_inp;
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1153_assgn1153);
    assign z4121_assgn4121 = dec_2_inp;
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1155_assgn1155);
    assign z4125_assgn4125 = dec_1_inp;
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1157_assgn1157);
    assign z4129_assgn4129 = dec_1_inp;
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1159_assgn1159);
    assign z4133_assgn4133 = dec_1_inp;
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1161_assgn1161);
    assign z4137_assgn4137 = dec_1_inp;
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1163_assgn1163);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign z4149_assgn4149 = dec_1_inp;
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << z1173_assgn1173);
    assign z4153_assgn4153 = dec_1_inp;
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << z1175_assgn1175);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (v_r1_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul3_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul3_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul3_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4173_assgn4173 = dec_2_inp;
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1193_assgn1193);
    assign z4177_assgn4177 = dec_2_inp;
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1195_assgn1195);
    assign z4181_assgn4181 = dec_1_inp;
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> z1197_assgn1197);
    assign z4185_assgn4185 = dec_1_inp;
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> z1199_assgn1199);
    assign z4189_assgn4189 = dec_1_inp;
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1201_assgn1201);
    assign z4193_assgn4193 = dec_1_inp;
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1203_assgn1203);
    assign z4197_assgn4197 = dec_2_inp;
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1205_assgn1205);
    assign z4201_assgn4201 = dec_2_inp;
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1207_assgn1207);
    assign z4205_assgn4205 = dec_1_inp;
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> z1209_assgn1209);
    assign z4209_assgn4209 = dec_1_inp;
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> z1211_assgn1211);
    assign z4213_assgn4213 = dec_1_inp;
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1213_assgn1213);
    assign z4217_assgn4217 = dec_1_inp;
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1215_assgn1215);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ d1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_hpc10_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4233_assgn4233 = r00_hpc10_G4_mul3_G16_inv0_G256_inv0;
    assign b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0 = (cxord_0_G4_mul3_G16_inv0_G256_inv0 ^ z1229_assgn1229);
    assign z4237_assgn4237 = r00_hpc10_G4_mul3_G16_inv0_G256_inv0;
    assign b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0 = (cxord_1_G4_mul3_G16_inv0_G256_inv0 ^ z1231_assgn1231);
    assign p2_hpc10_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4243_assgn4243 = r10_hpc10_G4_mul3_G16_inv0_G256_inv0;
    assign i1_hpc10_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc10_G4_mul3_G16_inv0_G256_inv0 ^ z1235_assgn1235);
    assign p3_hpc10_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4249_assgn4249 = r10_hpc10_G4_mul3_G16_inv0_G256_inv0;
    assign i2_hpc10_G4_mul3_G16_inv0_G256_inv0 = (p3_hpc10_G4_mul3_G16_inv0_G256_inv0 ^ z1239_assgn1239);
    assign p1_hpc10_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_hpc10_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (i1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (i2_hpc10_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_hpc10_G4_mul3_G16_inv0_G256_inv0_reg);
    assign r00_hpc11_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4265_assgn4265 = r00_hpc11_G4_mul3_G16_inv0_G256_inv0;
    assign b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ z1253_assgn1253);
    assign z4269_assgn4269 = r00_hpc11_G4_mul3_G16_inv0_G256_inv0;
    assign b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ z1255_assgn1255);
    assign p2_hpc11_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4275_assgn4275 = r10_hpc11_G4_mul3_G16_inv0_G256_inv0;
    assign i1_hpc11_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc11_G4_mul3_G16_inv0_G256_inv0 ^ z1259_assgn1259);
    assign p3_hpc11_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4281_assgn4281 = r10_hpc11_G4_mul3_G16_inv0_G256_inv0;
    assign i2_hpc11_G4_mul3_G16_inv0_G256_inv0 = (p3_hpc11_G4_mul3_G16_inv0_G256_inv0 ^ z1263_assgn1263);
    assign p1_hpc11_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_hpc11_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (i1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (i2_hpc11_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_hpc11_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_hpc12_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4301_assgn4301 = r00_hpc12_G4_mul3_G16_inv0_G256_inv0;
    assign b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0 = (d0_G4_mul3_G16_inv0_G256_inv0 ^ z1281_assgn1281);
    assign z4305_assgn4305 = r00_hpc12_G4_mul3_G16_inv0_G256_inv0;
    assign b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0 = (d1_G4_mul3_G16_inv0_G256_inv0 ^ z1283_assgn1283);
    assign p2_hpc12_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4311_assgn4311 = r10_hpc12_G4_mul3_G16_inv0_G256_inv0;
    assign i1_hpc12_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc12_G4_mul3_G16_inv0_G256_inv0 ^ z1287_assgn1287);
    assign p3_hpc12_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4317_assgn4317 = r10_hpc12_G4_mul3_G16_inv0_G256_inv0;
    assign i2_hpc12_G4_mul3_G16_inv0_G256_inv0 = (p3_hpc12_G4_mul3_G16_inv0_G256_inv0 ^ z1291_assgn1291);
    assign p1_hpc12_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0_reg & b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_hpc12_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0_reg & b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (i1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (i2_hpc12_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_hpc12_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z4333_assgn4333 = dec_1_inp;
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << z1305_assgn1305);
    assign z4337_assgn4337 = dec_1_inp;
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << z1307_assgn1307);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign z4345_assgn4345 = c0_G16_inv0_G256_inv0;
    assign c0xord0_G16_inv0_G256_inv0 = (z1314_assgn1314 ^ d0_G16_inv0_G256_inv0);
    assign z4349_assgn4349 = c1_G16_inv0_G256_inv0;
    assign c1xord1_G16_inv0_G256_inv0 = (z1316_assgn1316 ^ d1_G16_inv0_G256_inv0);
    assign z4353_assgn4353 = dec_2_inp;
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1317_assgn1317);
    assign z4357_assgn4357 = dec_2_inp;
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1319_assgn1319);
    assign z4361_assgn4361 = dec_1_inp;
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> z1321_assgn1321);
    assign z4365_assgn4365 = dec_1_inp;
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> z1323_assgn1323);
    assign z4369_assgn4369 = dec_1_inp;
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1325_assgn1325);
    assign z4373_assgn4373 = dec_1_inp;
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1327_assgn1327);
    assign z4377_assgn4377 = dec_1_inp;
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << z1329_assgn1329);
    assign z4381_assgn4381 = dec_1_inp;
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << z1331_assgn1331);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r60_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r70_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r80_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul4_G16_inv0_G256_inv0 = (r90_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul4_G16_inv0_G256_inv0 = (r100_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul4_G16_inv0_G256_inv0 = (r110_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4401_assgn4401 = dec_2_inp;
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1349_assgn1349);
    assign z4405_assgn4405 = dec_2_inp;
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1351_assgn1351);
    assign z4409_assgn4409 = dec_1_inp;
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> z1353_assgn1353);
    assign z4413_assgn4413 = dec_1_inp;
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> z1355_assgn1355);
    assign z4417_assgn4417 = dec_1_inp;
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1357_assgn1357);
    assign z4421_assgn4421 = dec_1_inp;
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1359_assgn1359);
    assign z4425_assgn4425 = dec_2_inp;
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1361_assgn1361);
    assign z4429_assgn4429 = dec_2_inp;
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1363_assgn1363);
    assign z4433_assgn4433 = dec_1_inp;
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> z1365_assgn1365);
    assign z4437_assgn4437 = dec_1_inp;
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> z1367_assgn1367);
    assign z4441_assgn4441 = dec_1_inp;
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1369_assgn1369);
    assign z4445_assgn4445 = dec_1_inp;
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1371_assgn1371);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ d1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_hpc10_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4461_assgn4461 = r00_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign b0_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0 = (cxord_0_G4_mul4_G16_inv0_G256_inv0 ^ z1385_assgn1385);
    assign z4465_assgn4465 = r00_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign b1_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0 = (cxord_1_G4_mul4_G16_inv0_G256_inv0 ^ z1387_assgn1387);
    assign z4469_assgn4469 = b1_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc10_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & z1389_assgn1389);
    assign z4473_assgn4473 = r10_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign i1_hpc10_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc10_G4_mul4_G16_inv0_G256_inv0 ^ z1391_assgn1391);
    assign z4477_assgn4477 = b0_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc10_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & z1393_assgn1393);
    assign z4481_assgn4481 = r10_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign i2_hpc10_G4_mul4_G16_inv0_G256_inv0 = (p3_hpc10_G4_mul4_G16_inv0_G256_inv0 ^ z1395_assgn1395);
    assign z4485_assgn4485 = b0_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc10_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & z1397_assgn1397);
    assign z4489_assgn4489 = b1_preshared_hpc10_G4_mul4_G16_inv0_G256_inv0;
    assign p4_hpc10_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & z1399_assgn1399);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (i1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (i2_hpc10_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_hpc10_G4_mul4_G16_inv0_G256_inv0_reg);
    assign r00_hpc11_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4501_assgn4501 = r00_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign b0_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ z1409_assgn1409);
    assign z4505_assgn4505 = r00_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign b1_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ z1411_assgn1411);
    assign z4509_assgn4509 = b1_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc11_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & z1413_assgn1413);
    assign z4513_assgn4513 = r10_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign i1_hpc11_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc11_G4_mul4_G16_inv0_G256_inv0 ^ z1415_assgn1415);
    assign z4517_assgn4517 = b0_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc11_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & z1417_assgn1417);
    assign z4521_assgn4521 = r10_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign i2_hpc11_G4_mul4_G16_inv0_G256_inv0 = (p3_hpc11_G4_mul4_G16_inv0_G256_inv0 ^ z1419_assgn1419);
    assign z4525_assgn4525 = b0_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc11_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & z1421_assgn1421);
    assign z4529_assgn4529 = b1_preshared_hpc11_G4_mul4_G16_inv0_G256_inv0;
    assign p4_hpc11_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & z1423_assgn1423);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (i1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (i2_hpc11_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_hpc11_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_hpc12_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4545_assgn4545 = r00_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign b0_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0 = (d0_G4_mul4_G16_inv0_G256_inv0 ^ z1437_assgn1437);
    assign z4549_assgn4549 = r00_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign b1_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0 = (d1_G4_mul4_G16_inv0_G256_inv0 ^ z1439_assgn1439);
    assign z4553_assgn4553 = b1_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc12_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & z1441_assgn1441);
    assign z4557_assgn4557 = r10_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign i1_hpc12_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc12_G4_mul4_G16_inv0_G256_inv0 ^ z1443_assgn1443);
    assign z4561_assgn4561 = b0_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc12_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & z1445_assgn1445);
    assign z4565_assgn4565 = r10_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign i2_hpc12_G4_mul4_G16_inv0_G256_inv0 = (p3_hpc12_G4_mul4_G16_inv0_G256_inv0 ^ z1447_assgn1447);
    assign z4569_assgn4569 = b0_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc12_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & z1449_assgn1449);
    assign z4573_assgn4573 = b1_preshared_hpc12_G4_mul4_G16_inv0_G256_inv0;
    assign p4_hpc12_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & z1451_assgn1451);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (i1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (i2_hpc12_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_hpc12_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z4585_assgn4585 = dec_1_inp;
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << z1461_assgn1461);
    assign z4589_assgn4589 = dec_1_inp;
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << z1463_assgn1463);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r120_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r130_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r140_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul5_G16_inv0_G256_inv0 = (r150_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul5_G16_inv0_G256_inv0 = (r160_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul5_G16_inv0_G256_inv0 = (r170_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4609_assgn4609 = dec_2_inp;
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1481_assgn1481);
    assign z4613_assgn4613 = dec_2_inp;
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1483_assgn1483);
    assign z4617_assgn4617 = dec_1_inp;
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> z1485_assgn1485);
    assign z4621_assgn4621 = dec_1_inp;
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> z1487_assgn1487);
    assign z4625_assgn4625 = dec_1_inp;
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1489_assgn1489);
    assign z4629_assgn4629 = dec_1_inp;
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1491_assgn1491);
    assign z4633_assgn4633 = dec_2_inp;
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1493_assgn1493);
    assign z4637_assgn4637 = dec_2_inp;
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1495_assgn1495);
    assign z4641_assgn4641 = dec_1_inp;
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> z1497_assgn1497);
    assign z4645_assgn4645 = dec_1_inp;
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> z1499_assgn1499);
    assign z4649_assgn4649 = dec_1_inp;
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1501_assgn1501);
    assign z4653_assgn4653 = dec_1_inp;
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1503_assgn1503);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ d1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_hpc10_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4669_assgn4669 = r00_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign b0_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0 = (cxord_0_G4_mul5_G16_inv0_G256_inv0 ^ z1517_assgn1517);
    assign z4673_assgn4673 = r00_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign b1_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0 = (cxord_1_G4_mul5_G16_inv0_G256_inv0 ^ z1519_assgn1519);
    assign z4677_assgn4677 = b1_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc10_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & z1521_assgn1521);
    assign z4681_assgn4681 = r10_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign i1_hpc10_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc10_G4_mul5_G16_inv0_G256_inv0 ^ z1523_assgn1523);
    assign z4685_assgn4685 = b0_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc10_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & z1525_assgn1525);
    assign z4689_assgn4689 = r10_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign i2_hpc10_G4_mul5_G16_inv0_G256_inv0 = (p3_hpc10_G4_mul5_G16_inv0_G256_inv0 ^ z1527_assgn1527);
    assign z4693_assgn4693 = b0_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc10_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & z1529_assgn1529);
    assign z4697_assgn4697 = b1_preshared_hpc10_G4_mul5_G16_inv0_G256_inv0;
    assign p4_hpc10_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & z1531_assgn1531);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (i1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (i2_hpc10_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_hpc10_G4_mul5_G16_inv0_G256_inv0_reg);
    assign r00_hpc11_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4709_assgn4709 = r00_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign b0_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ z1541_assgn1541);
    assign z4713_assgn4713 = r00_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign b1_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ z1543_assgn1543);
    assign z4717_assgn4717 = b1_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc11_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & z1545_assgn1545);
    assign z4721_assgn4721 = r10_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign i1_hpc11_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc11_G4_mul5_G16_inv0_G256_inv0 ^ z1547_assgn1547);
    assign z4725_assgn4725 = b0_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc11_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & z1549_assgn1549);
    assign z4729_assgn4729 = r10_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign i2_hpc11_G4_mul5_G16_inv0_G256_inv0 = (p3_hpc11_G4_mul5_G16_inv0_G256_inv0 ^ z1551_assgn1551);
    assign z4733_assgn4733 = b0_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc11_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & z1553_assgn1553);
    assign z4737_assgn4737 = b1_preshared_hpc11_G4_mul5_G16_inv0_G256_inv0;
    assign p4_hpc11_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & z1555_assgn1555);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (i1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (i2_hpc11_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_hpc11_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_hpc12_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign z4753_assgn4753 = r00_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign b0_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0 = (d0_G4_mul5_G16_inv0_G256_inv0 ^ z1569_assgn1569);
    assign z4757_assgn4757 = r00_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign b1_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0 = (d1_G4_mul5_G16_inv0_G256_inv0 ^ z1571_assgn1571);
    assign z4761_assgn4761 = b1_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc12_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & z1573_assgn1573);
    assign z4765_assgn4765 = r10_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign i1_hpc12_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc12_G4_mul5_G16_inv0_G256_inv0 ^ z1575_assgn1575);
    assign z4769_assgn4769 = b0_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc12_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & z1577_assgn1577);
    assign z4773_assgn4773 = r10_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign i2_hpc12_G4_mul5_G16_inv0_G256_inv0 = (p3_hpc12_G4_mul5_G16_inv0_G256_inv0 ^ z1579_assgn1579);
    assign z4777_assgn4777 = b0_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc12_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & z1581_assgn1581);
    assign z4781_assgn4781 = b1_preshared_hpc12_G4_mul5_G16_inv0_G256_inv0;
    assign p4_hpc12_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & z1583_assgn1583);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (i1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (i2_hpc12_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_hpc12_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z4793_assgn4793 = dec_1_inp;
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << z1593_assgn1593);
    assign z4797_assgn4797 = dec_1_inp;
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << z1595_assgn1595);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign z4805_assgn4805 = dec_2_inp;
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << z1601_assgn1601);
    assign z4809_assgn4809 = dec_2_inp;
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << z1603_assgn1603);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign r00_G16_mul1_G256_inv0 = (r36_inp % dec_16_inp);
    assign v_r1_G16_mul1_G256_inv0 = (r37_inp % dec_16_inp);
    assign r20_G16_mul1_G256_inv0 = (r38_inp % dec_16_inp);
    assign r30_G16_mul1_G256_inv0 = (r39_inp % dec_16_inp);
    assign r40_G16_mul1_G256_inv0 = (r40_inp % dec_16_inp);
    assign r50_G16_mul1_G256_inv0 = (r41_inp % dec_16_inp);
    assign r60_G16_mul1_G256_inv0 = (r42_inp % dec_16_inp);
    assign r70_G16_mul1_G256_inv0 = (r43_inp % dec_16_inp);
    assign r80_G16_mul1_G256_inv0 = (r44_inp % dec_16_inp);
    assign r90_G16_mul1_G256_inv0 = (r45_inp % dec_16_inp);
    assign r100_G16_mul1_G256_inv0 = (r46_inp % dec_16_inp);
    assign r110_G16_mul1_G256_inv0 = (r47_inp % dec_16_inp);
    assign r120_G16_mul1_G256_inv0 = (r48_inp % dec_16_inp);
    assign r130_G16_mul1_G256_inv0 = (r49_inp % dec_16_inp);
    assign r140_G16_mul1_G256_inv0 = (r50_inp % dec_16_inp);
    assign r150_G16_mul1_G256_inv0 = (r51_inp % dec_16_inp);
    assign r160_G16_mul1_G256_inv0 = (r52_inp % dec_16_inp);
    assign r170_G16_mul1_G256_inv0 = (r53_inp % dec_16_inp);
    assign z4853_assgn4853 = dec_12_inp;
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1645_assgn1645);
    assign z4857_assgn4857 = dec_12_inp;
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1647_assgn1647);
    assign z4861_assgn4861 = dec_2_inp;
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> z1649_assgn1649);
    assign z4865_assgn4865 = dec_2_inp;
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> z1651_assgn1651);
    assign z4869_assgn4869 = dec_3_inp;
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1653_assgn1653);
    assign z4873_assgn4873 = dec_3_inp;
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1655_assgn1655);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (v_r1_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign z4909_assgn4909 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1689_assgn1689);
    assign z4913_assgn4913 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1691_assgn1691);
    assign z4917_assgn4917 = dec_1_inp;
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> z1693_assgn1693);
    assign z4921_assgn4921 = dec_1_inp;
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> z1695_assgn1695);
    assign z4925_assgn4925 = dec_1_inp;
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1697_assgn1697);
    assign z4929_assgn4929 = dec_1_inp;
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1699_assgn1699);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ d1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_hpc10_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul1_G256_inv0);
    assign b1_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul1_G256_inv0);
    assign z4961_assgn4961 = b1_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc10_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1729_assgn1729);
    assign z4965_assgn4965 = r10_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign i1_hpc10_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc10_G4_mul0_G16_mul1_G256_inv0 ^ z1731_assgn1731);
    assign z4969_assgn4969 = b0_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc10_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1733_assgn1733);
    assign z4973_assgn4973 = r10_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign i2_hpc10_G4_mul0_G16_mul1_G256_inv0 = (p3_hpc10_G4_mul0_G16_mul1_G256_inv0 ^ z1735_assgn1735);
    assign z4977_assgn4977 = b0_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc10_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1737_assgn1737);
    assign z4981_assgn4981 = b1_preshared_hpc10_G4_mul0_G16_mul1_G256_inv0;
    assign p4_hpc10_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1739_assgn1739);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (i1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (i2_hpc10_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_hpc10_G4_mul0_G16_mul1_G256_inv0_reg);
    assign r00_hpc11_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul1_G256_inv0);
    assign b1_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul1_G256_inv0);
    assign z4997_assgn4997 = b1_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc11_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1753_assgn1753);
    assign z5001_assgn5001 = r10_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign i1_hpc11_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc11_G4_mul0_G16_mul1_G256_inv0 ^ z1755_assgn1755);
    assign z5005_assgn5005 = b0_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc11_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1757_assgn1757);
    assign z5009_assgn5009 = r10_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign i2_hpc11_G4_mul0_G16_mul1_G256_inv0 = (p3_hpc11_G4_mul0_G16_mul1_G256_inv0 ^ z1759_assgn1759);
    assign z5013_assgn5013 = b0_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc11_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1761_assgn1761);
    assign z5017_assgn5017 = b1_preshared_hpc11_G4_mul0_G16_mul1_G256_inv0;
    assign p4_hpc11_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1763_assgn1763);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (i1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (i2_hpc11_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_hpc11_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_hpc12_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0 = (d0_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul1_G256_inv0);
    assign b1_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0 = (d1_G4_mul0_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul1_G256_inv0);
    assign z5037_assgn5037 = b1_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc12_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1781_assgn1781);
    assign z5041_assgn5041 = r10_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign i1_hpc12_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc12_G4_mul0_G16_mul1_G256_inv0 ^ z1783_assgn1783);
    assign z5045_assgn5045 = b0_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc12_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1785_assgn1785);
    assign z5049_assgn5049 = r10_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign i2_hpc12_G4_mul0_G16_mul1_G256_inv0 = (p3_hpc12_G4_mul0_G16_mul1_G256_inv0 ^ z1787_assgn1787);
    assign z5053_assgn5053 = b0_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc12_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1789_assgn1789);
    assign z5057_assgn5057 = b1_preshared_hpc12_G4_mul0_G16_mul1_G256_inv0;
    assign p4_hpc12_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1791_assgn1791);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (i1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (i2_hpc12_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_hpc12_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z5069_assgn5069 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << z1801_assgn1801);
    assign z5073_assgn5073 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << z1803_assgn1803);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign z5081_assgn5081 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1809_assgn1809);
    assign z5085_assgn5085 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1811_assgn1811);
    assign z5089_assgn5089 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1813_assgn1813);
    assign z5093_assgn5093 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1815_assgn1815);
    assign z5097_assgn5097 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1817_assgn1817);
    assign z5101_assgn5101 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1819_assgn1819);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z5113_assgn5113 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << z1829_assgn1829);
    assign z5117_assgn5117 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << z1831_assgn1831);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r60_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r70_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r80_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul1_G256_inv0 = (r90_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul1_G256_inv0 = (r100_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul1_G256_inv0 = (r110_G16_mul1_G256_inv0 % dec_4_inp);
    assign z5137_assgn5137 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1849_assgn1849);
    assign z5141_assgn5141 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1851_assgn1851);
    assign z5145_assgn5145 = dec_1_inp;
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> z1853_assgn1853);
    assign z5149_assgn5149 = dec_1_inp;
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> z1855_assgn1855);
    assign z5153_assgn5153 = dec_1_inp;
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1857_assgn1857);
    assign z5157_assgn5157 = dec_1_inp;
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1859_assgn1859);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ d1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_hpc10_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0 = (cxord_0_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul1_G256_inv0);
    assign b1_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0 = (cxord_1_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul1_G256_inv0);
    assign z5189_assgn5189 = b1_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc10_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1889_assgn1889);
    assign z5193_assgn5193 = r10_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign i1_hpc10_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc10_G4_mul1_G16_mul1_G256_inv0 ^ z1891_assgn1891);
    assign z5197_assgn5197 = b0_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc10_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1893_assgn1893);
    assign z5201_assgn5201 = r10_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign i2_hpc10_G4_mul1_G16_mul1_G256_inv0 = (p3_hpc10_G4_mul1_G16_mul1_G256_inv0 ^ z1895_assgn1895);
    assign z5205_assgn5205 = b0_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc10_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1897_assgn1897);
    assign z5209_assgn5209 = b1_preshared_hpc10_G4_mul1_G16_mul1_G256_inv0;
    assign p4_hpc10_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1899_assgn1899);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (i1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (i2_hpc10_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_hpc10_G4_mul1_G16_mul1_G256_inv0_reg);
    assign r00_hpc11_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul1_G256_inv0);
    assign b1_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul1_G256_inv0);
    assign z5225_assgn5225 = b1_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc11_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1913_assgn1913);
    assign z5229_assgn5229 = r10_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign i1_hpc11_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc11_G4_mul1_G16_mul1_G256_inv0 ^ z1915_assgn1915);
    assign z5233_assgn5233 = b0_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc11_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1917_assgn1917);
    assign z5237_assgn5237 = r10_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign i2_hpc11_G4_mul1_G16_mul1_G256_inv0 = (p3_hpc11_G4_mul1_G16_mul1_G256_inv0 ^ z1919_assgn1919);
    assign z5241_assgn5241 = b0_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc11_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1921_assgn1921);
    assign z5245_assgn5245 = b1_preshared_hpc11_G4_mul1_G16_mul1_G256_inv0;
    assign p4_hpc11_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1923_assgn1923);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (i1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (i2_hpc11_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_hpc11_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_hpc12_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0 = (d0_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul1_G256_inv0);
    assign b1_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0 = (d1_G4_mul1_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul1_G256_inv0);
    assign z5265_assgn5265 = b1_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc12_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1941_assgn1941);
    assign z5269_assgn5269 = r10_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign i1_hpc12_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc12_G4_mul1_G16_mul1_G256_inv0 ^ z1943_assgn1943);
    assign z5273_assgn5273 = b0_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc12_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1945_assgn1945);
    assign z5277_assgn5277 = r10_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign i2_hpc12_G4_mul1_G16_mul1_G256_inv0 = (p3_hpc12_G4_mul1_G16_mul1_G256_inv0 ^ z1947_assgn1947);
    assign z5281_assgn5281 = b0_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc12_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1949_assgn1949);
    assign z5285_assgn5285 = b1_preshared_hpc12_G4_mul1_G16_mul1_G256_inv0;
    assign p4_hpc12_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1951_assgn1951);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (i1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (i2_hpc12_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_hpc12_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z5297_assgn5297 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << z1961_assgn1961);
    assign z5301_assgn5301 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << z1963_assgn1963);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r120_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r130_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r140_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul1_G256_inv0 = (r150_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul1_G256_inv0 = (r160_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul1_G256_inv0 = (r170_G16_mul1_G256_inv0 % dec_4_inp);
    assign z5325_assgn5325 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1985_assgn1985);
    assign z5329_assgn5329 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1987_assgn1987);
    assign z5333_assgn5333 = dec_1_inp;
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> z1989_assgn1989);
    assign z5337_assgn5337 = dec_1_inp;
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> z1991_assgn1991);
    assign z5341_assgn5341 = dec_1_inp;
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1993_assgn1993);
    assign z5345_assgn5345 = dec_1_inp;
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1995_assgn1995);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ d1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_hpc10_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0 = (cxord_0_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul1_G256_inv0);
    assign b1_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0 = (cxord_1_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul1_G256_inv0);
    assign z5377_assgn5377 = b1_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc10_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z2025_assgn2025);
    assign z5381_assgn5381 = r10_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign i1_hpc10_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc10_G4_mul2_G16_mul1_G256_inv0 ^ z2027_assgn2027);
    assign z5385_assgn5385 = b0_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc10_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z2029_assgn2029);
    assign z5389_assgn5389 = r10_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign i2_hpc10_G4_mul2_G16_mul1_G256_inv0 = (p3_hpc10_G4_mul2_G16_mul1_G256_inv0 ^ z2031_assgn2031);
    assign z5393_assgn5393 = b0_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc10_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z2033_assgn2033);
    assign z5397_assgn5397 = b1_preshared_hpc10_G4_mul2_G16_mul1_G256_inv0;
    assign p4_hpc10_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z2035_assgn2035);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (i1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (i2_hpc10_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_hpc10_G4_mul2_G16_mul1_G256_inv0_reg);
    assign r00_hpc11_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul1_G256_inv0);
    assign b1_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul1_G256_inv0);
    assign z5413_assgn5413 = b1_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc11_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z2049_assgn2049);
    assign z5417_assgn5417 = r10_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign i1_hpc11_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc11_G4_mul2_G16_mul1_G256_inv0 ^ z2051_assgn2051);
    assign z5421_assgn5421 = b0_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc11_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z2053_assgn2053);
    assign z5425_assgn5425 = r10_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign i2_hpc11_G4_mul2_G16_mul1_G256_inv0 = (p3_hpc11_G4_mul2_G16_mul1_G256_inv0 ^ z2055_assgn2055);
    assign z5429_assgn5429 = b0_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc11_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z2057_assgn2057);
    assign z5433_assgn5433 = b1_preshared_hpc11_G4_mul2_G16_mul1_G256_inv0;
    assign p4_hpc11_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z2059_assgn2059);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (i1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (i2_hpc11_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_hpc11_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_hpc12_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0 = (d0_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul1_G256_inv0);
    assign b1_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0 = (d1_G4_mul2_G16_mul1_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul1_G256_inv0);
    assign z5453_assgn5453 = b1_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc12_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z2077_assgn2077);
    assign z5457_assgn5457 = r10_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign i1_hpc12_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc12_G4_mul2_G16_mul1_G256_inv0 ^ z2079_assgn2079);
    assign z5461_assgn5461 = b0_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc12_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z2081_assgn2081);
    assign z5465_assgn5465 = r10_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign i2_hpc12_G4_mul2_G16_mul1_G256_inv0 = (p3_hpc12_G4_mul2_G16_mul1_G256_inv0 ^ z2083_assgn2083);
    assign z5469_assgn5469 = b0_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc12_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z2085_assgn2085);
    assign z5473_assgn5473 = b1_preshared_hpc12_G4_mul2_G16_mul1_G256_inv0;
    assign p4_hpc12_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z2087_assgn2087);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (i1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (i2_hpc12_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_hpc12_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z5485_assgn5485 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << z2097_assgn2097);
    assign z5489_assgn5489 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << z2099_assgn2099);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign z5501_assgn5501 = dec_2_inp;
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << z2109_assgn2109);
    assign z5505_assgn5505 = dec_2_inp;
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << z2111_assgn2111);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign r00_G16_mul2_G256_inv0 = (r54_inp % dec_16_inp);
    assign v_r1_G16_mul2_G256_inv0 = (r55_inp % dec_16_inp);
    assign r20_G16_mul2_G256_inv0 = (r56_inp % dec_16_inp);
    assign r30_G16_mul2_G256_inv0 = (r57_inp % dec_16_inp);
    assign r40_G16_mul2_G256_inv0 = (r58_inp % dec_16_inp);
    assign r50_G16_mul2_G256_inv0 = (r59_inp % dec_16_inp);
    assign r60_G16_mul2_G256_inv0 = (r60_inp % dec_16_inp);
    assign r70_G16_mul2_G256_inv0 = (r61_inp % dec_16_inp);
    assign r80_G16_mul2_G256_inv0 = (r62_inp % dec_16_inp);
    assign r90_G16_mul2_G256_inv0 = (r63_inp % dec_16_inp);
    assign r100_G16_mul2_G256_inv0 = (r64_inp % dec_16_inp);
    assign r110_G16_mul2_G256_inv0 = (r65_inp % dec_16_inp);
    assign r120_G16_mul2_G256_inv0 = (r66_inp % dec_16_inp);
    assign r130_G16_mul2_G256_inv0 = (r67_inp % dec_16_inp);
    assign r140_G16_mul2_G256_inv0 = (r68_inp % dec_16_inp);
    assign r150_G16_mul2_G256_inv0 = (r69_inp % dec_16_inp);
    assign r160_G16_mul2_G256_inv0 = (r70_inp % dec_16_inp);
    assign r170_G16_mul2_G256_inv0 = (r71_inp % dec_16_inp);
    assign z5549_assgn5549 = dec_12_inp;
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2153_assgn2153);
    assign z5553_assgn5553 = dec_12_inp;
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2155_assgn2155);
    assign z5557_assgn5557 = dec_2_inp;
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> z2157_assgn2157);
    assign z5561_assgn5561 = dec_2_inp;
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> z2159_assgn2159);
    assign z5565_assgn5565 = dec_3_inp;
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2161_assgn2161);
    assign z5569_assgn5569 = dec_3_inp;
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2163_assgn2163);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (v_r1_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign z5605_assgn5605 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2197_assgn2197);
    assign z5609_assgn5609 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2199_assgn2199);
    assign z5613_assgn5613 = dec_1_inp;
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> z2201_assgn2201);
    assign z5617_assgn5617 = dec_1_inp;
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> z2203_assgn2203);
    assign z5621_assgn5621 = dec_1_inp;
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2205_assgn2205);
    assign z5625_assgn5625 = dec_1_inp;
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2207_assgn2207);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ d1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_hpc10_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul2_G256_inv0);
    assign b1_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul0_G16_mul2_G256_inv0);
    assign z5657_assgn5657 = b1_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc10_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z2237_assgn2237);
    assign z5661_assgn5661 = r10_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign i1_hpc10_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc10_G4_mul0_G16_mul2_G256_inv0 ^ z2239_assgn2239);
    assign z5665_assgn5665 = b0_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc10_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z2241_assgn2241);
    assign z5669_assgn5669 = r10_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign i2_hpc10_G4_mul0_G16_mul2_G256_inv0 = (p3_hpc10_G4_mul0_G16_mul2_G256_inv0 ^ z2243_assgn2243);
    assign z5673_assgn5673 = b0_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc10_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z2245_assgn2245);
    assign z5677_assgn5677 = b1_preshared_hpc10_G4_mul0_G16_mul2_G256_inv0;
    assign p4_hpc10_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z2247_assgn2247);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (i1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (i2_hpc10_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_hpc10_G4_mul0_G16_mul2_G256_inv0_reg);
    assign r00_hpc11_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul2_G256_inv0);
    assign b1_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul0_G16_mul2_G256_inv0);
    assign z5693_assgn5693 = b1_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc11_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z2261_assgn2261);
    assign z5697_assgn5697 = r10_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign i1_hpc11_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc11_G4_mul0_G16_mul2_G256_inv0 ^ z2263_assgn2263);
    assign z5701_assgn5701 = b0_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc11_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z2265_assgn2265);
    assign z5705_assgn5705 = r10_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign i2_hpc11_G4_mul0_G16_mul2_G256_inv0 = (p3_hpc11_G4_mul0_G16_mul2_G256_inv0 ^ z2267_assgn2267);
    assign z5709_assgn5709 = b0_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc11_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z2269_assgn2269);
    assign z5713_assgn5713 = b1_preshared_hpc11_G4_mul0_G16_mul2_G256_inv0;
    assign p4_hpc11_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z2271_assgn2271);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (i1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (i2_hpc11_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_hpc11_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_hpc12_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0 = (d0_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul2_G256_inv0);
    assign b1_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0 = (d1_G4_mul0_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul0_G16_mul2_G256_inv0);
    assign z5733_assgn5733 = b1_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc12_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z2289_assgn2289);
    assign z5737_assgn5737 = r10_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign i1_hpc12_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc12_G4_mul0_G16_mul2_G256_inv0 ^ z2291_assgn2291);
    assign z5741_assgn5741 = b0_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc12_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z2293_assgn2293);
    assign z5745_assgn5745 = r10_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign i2_hpc12_G4_mul0_G16_mul2_G256_inv0 = (p3_hpc12_G4_mul0_G16_mul2_G256_inv0 ^ z2295_assgn2295);
    assign z5749_assgn5749 = b0_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc12_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z2297_assgn2297);
    assign z5753_assgn5753 = b1_preshared_hpc12_G4_mul0_G16_mul2_G256_inv0;
    assign p4_hpc12_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z2299_assgn2299);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (i1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (i2_hpc12_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_hpc12_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z5765_assgn5765 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << z2309_assgn2309);
    assign z5769_assgn5769 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << z2311_assgn2311);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign z5777_assgn5777 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2317_assgn2317);
    assign z5781_assgn5781 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2319_assgn2319);
    assign z5785_assgn5785 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2321_assgn2321);
    assign z5789_assgn5789 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2323_assgn2323);
    assign z5793_assgn5793 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2325_assgn2325);
    assign z5797_assgn5797 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2327_assgn2327);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z5809_assgn5809 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << z2337_assgn2337);
    assign z5813_assgn5813 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << z2339_assgn2339);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r60_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r70_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r80_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul2_G256_inv0 = (r90_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul2_G256_inv0 = (r100_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul2_G256_inv0 = (r110_G16_mul2_G256_inv0 % dec_4_inp);
    assign z5833_assgn5833 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2357_assgn2357);
    assign z5837_assgn5837 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2359_assgn2359);
    assign z5841_assgn5841 = dec_1_inp;
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> z2361_assgn2361);
    assign z5845_assgn5845 = dec_1_inp;
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> z2363_assgn2363);
    assign z5849_assgn5849 = dec_1_inp;
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2365_assgn2365);
    assign z5853_assgn5853 = dec_1_inp;
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2367_assgn2367);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ d1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_hpc10_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0 = (cxord_0_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul2_G256_inv0);
    assign b1_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0 = (cxord_1_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul1_G16_mul2_G256_inv0);
    assign z5885_assgn5885 = b1_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc10_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2397_assgn2397);
    assign z5889_assgn5889 = r10_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign i1_hpc10_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc10_G4_mul1_G16_mul2_G256_inv0 ^ z2399_assgn2399);
    assign z5893_assgn5893 = b0_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc10_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2401_assgn2401);
    assign z5897_assgn5897 = r10_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign i2_hpc10_G4_mul1_G16_mul2_G256_inv0 = (p3_hpc10_G4_mul1_G16_mul2_G256_inv0 ^ z2403_assgn2403);
    assign z5901_assgn5901 = b0_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc10_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2405_assgn2405);
    assign z5905_assgn5905 = b1_preshared_hpc10_G4_mul1_G16_mul2_G256_inv0;
    assign p4_hpc10_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2407_assgn2407);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (i1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (i2_hpc10_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_hpc10_G4_mul1_G16_mul2_G256_inv0_reg);
    assign r00_hpc11_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul2_G256_inv0);
    assign b1_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul1_G16_mul2_G256_inv0);
    assign z5921_assgn5921 = b1_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc11_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2421_assgn2421);
    assign z5925_assgn5925 = r10_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign i1_hpc11_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc11_G4_mul1_G16_mul2_G256_inv0 ^ z2423_assgn2423);
    assign z5929_assgn5929 = b0_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc11_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2425_assgn2425);
    assign z5933_assgn5933 = r10_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign i2_hpc11_G4_mul1_G16_mul2_G256_inv0 = (p3_hpc11_G4_mul1_G16_mul2_G256_inv0 ^ z2427_assgn2427);
    assign z5937_assgn5937 = b0_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc11_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2429_assgn2429);
    assign z5941_assgn5941 = b1_preshared_hpc11_G4_mul1_G16_mul2_G256_inv0;
    assign p4_hpc11_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2431_assgn2431);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (i1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (i2_hpc11_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_hpc11_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_hpc12_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0 = (d0_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul2_G256_inv0);
    assign b1_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0 = (d1_G4_mul1_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul1_G16_mul2_G256_inv0);
    assign z5961_assgn5961 = b1_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc12_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2449_assgn2449);
    assign z5965_assgn5965 = r10_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign i1_hpc12_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc12_G4_mul1_G16_mul2_G256_inv0 ^ z2451_assgn2451);
    assign z5969_assgn5969 = b0_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc12_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2453_assgn2453);
    assign z5973_assgn5973 = r10_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign i2_hpc12_G4_mul1_G16_mul2_G256_inv0 = (p3_hpc12_G4_mul1_G16_mul2_G256_inv0 ^ z2455_assgn2455);
    assign z5977_assgn5977 = b0_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc12_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2457_assgn2457);
    assign z5981_assgn5981 = b1_preshared_hpc12_G4_mul1_G16_mul2_G256_inv0;
    assign p4_hpc12_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2459_assgn2459);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (i1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (i2_hpc12_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_hpc12_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z5993_assgn5993 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << z2469_assgn2469);
    assign z5997_assgn5997 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << z2471_assgn2471);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r120_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r130_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r140_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul2_G256_inv0 = (r150_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul2_G256_inv0 = (r160_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul2_G256_inv0 = (r170_G16_mul2_G256_inv0 % dec_4_inp);
    assign z6021_assgn6021 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2493_assgn2493);
    assign z6025_assgn6025 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2495_assgn2495);
    assign z6029_assgn6029 = dec_1_inp;
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> z2497_assgn2497);
    assign z6033_assgn6033 = dec_1_inp;
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> z2499_assgn2499);
    assign z6037_assgn6037 = dec_1_inp;
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2501_assgn2501);
    assign z6041_assgn6041 = dec_1_inp;
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2503_assgn2503);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ d1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_hpc10_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc10_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0 = (cxord_0_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul2_G256_inv0);
    assign b1_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0 = (cxord_1_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc10_G4_mul2_G16_mul2_G256_inv0);
    assign z6073_assgn6073 = b1_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc10_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2533_assgn2533);
    assign z6077_assgn6077 = r10_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign i1_hpc10_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc10_G4_mul2_G16_mul2_G256_inv0 ^ z2535_assgn2535);
    assign z6081_assgn6081 = b0_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc10_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2537_assgn2537);
    assign z6085_assgn6085 = r10_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign i2_hpc10_G4_mul2_G16_mul2_G256_inv0 = (p3_hpc10_G4_mul2_G16_mul2_G256_inv0 ^ z2539_assgn2539);
    assign z6089_assgn6089 = b0_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc10_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2541_assgn2541);
    assign z6093_assgn6093 = b1_preshared_hpc10_G4_mul2_G16_mul2_G256_inv0;
    assign p4_hpc10_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2543_assgn2543);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (i1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (i2_hpc10_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_hpc10_G4_mul2_G16_mul2_G256_inv0_reg);
    assign r00_hpc11_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc11_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul2_G256_inv0);
    assign b1_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc11_G4_mul2_G16_mul2_G256_inv0);
    assign z6109_assgn6109 = b1_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc11_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2557_assgn2557);
    assign z6113_assgn6113 = r10_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign i1_hpc11_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc11_G4_mul2_G16_mul2_G256_inv0 ^ z2559_assgn2559);
    assign z6117_assgn6117 = b0_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc11_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2561_assgn2561);
    assign z6121_assgn6121 = r10_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign i2_hpc11_G4_mul2_G16_mul2_G256_inv0 = (p3_hpc11_G4_mul2_G16_mul2_G256_inv0 ^ z2563_assgn2563);
    assign z6125_assgn6125 = b0_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc11_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2565_assgn2565);
    assign z6129_assgn6129 = b1_preshared_hpc11_G4_mul2_G16_mul2_G256_inv0;
    assign p4_hpc11_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2567_assgn2567);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (i1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (i2_hpc11_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_hpc11_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_hpc12_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_hpc12_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign b0_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0 = (d0_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul2_G256_inv0);
    assign b1_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0 = (d1_G4_mul2_G16_mul2_G256_inv0 ^ r00_hpc12_G4_mul2_G16_mul2_G256_inv0);
    assign z6149_assgn6149 = b1_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc12_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2585_assgn2585);
    assign z6153_assgn6153 = r10_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign i1_hpc12_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc12_G4_mul2_G16_mul2_G256_inv0 ^ z2587_assgn2587);
    assign z6157_assgn6157 = b0_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc12_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2589_assgn2589);
    assign z6161_assgn6161 = r10_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign i2_hpc12_G4_mul2_G16_mul2_G256_inv0 = (p3_hpc12_G4_mul2_G16_mul2_G256_inv0 ^ z2591_assgn2591);
    assign z6165_assgn6165 = b0_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc12_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2593_assgn2593);
    assign z6169_assgn6169 = b1_preshared_hpc12_G4_mul2_G16_mul2_G256_inv0;
    assign p4_hpc12_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2595_assgn2595);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (i1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (i2_hpc12_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_hpc12_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z6181_assgn6181 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << z2605_assgn2605);
    assign z6185_assgn6185 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << z2607_assgn2607);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign z6197_assgn6197 = dec_2_inp;
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << z2617_assgn2617);
    assign z6201_assgn6201 = dec_2_inp;
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << z2619_assgn2619);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign z6209_assgn6209 = dec_4_inp;
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << z2625_assgn2625);
    assign z6213_assgn6213 = dec_4_inp;
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << z2627_assgn2627);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign z6225_assgn6225 = dec_1_inp;
    assign cond1_G256_newbasis1 = (t4 & z2637_assgn2637);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign z6233_assgn6233 = yxorb1_G256_newbasis1;
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * z2643_assgn2643);
    assign z6237_assgn6237 = tempy1_G256_newbasis1;
    assign tempyIntoNegCond1_G256_newbasis1 = (z2646_assgn2646 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1);
    assign z6243_assgn6243 = dec_1_inp;
    assign x1_G256_newbasis1 = (t4 >> z2649_assgn2649);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign z6249_assgn6249 = dec_1_inp;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & z2653_assgn2653);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign z6255_assgn6255 = dec_3_inp;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ z2657_assgn2657);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempyIntoNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1);
    assign z6265_assgn6265 = dec_1_inp;
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> z2665_assgn2665);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign z6271_assgn6271 = dec_1_inp;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & z2669_assgn2669);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign z6277_assgn6277 = dec_4_inp;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ z2673_assgn2673);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempyIntoNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1);
    assign z6287_assgn6287 = dec_1_inp;
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> z2681_assgn2681);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign z6293_assgn6293 = dec_1_inp;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & z2685_assgn2685);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign z6299_assgn6299 = dec_220_inp;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ z2689_assgn2689);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempyIntoNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1);
    assign z6309_assgn6309 = dec_1_inp;
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> z2697_assgn2697);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign z6315_assgn6315 = dec_1_inp;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & z2701_assgn2701);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign z6321_assgn6321 = dec_11_inp;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ z2705_assgn2705);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempyIntoNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1);
    assign z6331_assgn6331 = dec_1_inp;
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> z2713_assgn2713);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign z6337_assgn6337 = dec_1_inp;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & z2717_assgn2717);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign z6343_assgn6343 = dec_158_inp;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ z2721_assgn2721);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempyIntoNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1);
    assign z6353_assgn6353 = dec_1_inp;
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> z2729_assgn2729);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign z6359_assgn6359 = dec_1_inp;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & z2733_assgn2733);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign z6365_assgn6365 = dec_45_inp;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ z2737_assgn2737);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempyIntoNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1);
    assign z6375_assgn6375 = dec_1_inp;
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> z2745_assgn2745);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign z6381_assgn6381 = dec_1_inp;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & z2749_assgn2749);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign z6387_assgn6387 = dec_88_inp;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ z2753_assgn2753);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempyIntoNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1);
    assign z6397_assgn6397 = dec_1_inp;
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> z2761_assgn2761);
    assign t6 = y8_G256_newbasis1;
    assign z_y_G256_newbasis1 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z6407_assgn6407 = dec_1_inp;
    assign z_cond1_G256_newbasis1 = (t5 & z2769_assgn2769);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z6415_assgn6415 = z_yxorb1_G256_newbasis1;
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z2775_assgn2775);
    assign z6419_assgn6419 = z_tempy1_G256_newbasis1;
    assign z_tempyIntoNegCond1_G256_newbasis1 = (z2778_assgn2778 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempyIntoNegCond1_G256_newbasis1);
    assign z6425_assgn6425 = dec_1_inp;
    assign z_x1_G256_newbasis1 = (t5 >> z2781_assgn2781);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z6431_assgn6431 = dec_1_inp;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & z2785_assgn2785);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z6437_assgn6437 = dec_3_inp;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ z2789_assgn2789);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempyIntoNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempyIntoNegCond2_G256_newbasis1);
    assign z6447_assgn6447 = dec_1_inp;
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> z2797_assgn2797);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z6453_assgn6453 = dec_1_inp;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & z2801_assgn2801);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z6459_assgn6459 = dec_4_inp;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ z2805_assgn2805);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempyIntoNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempyIntoNegCond3_G256_newbasis1);
    assign z6469_assgn6469 = dec_1_inp;
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> z2813_assgn2813);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z6475_assgn6475 = dec_1_inp;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & z2817_assgn2817);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z6481_assgn6481 = dec_220_inp;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ z2821_assgn2821);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempyIntoNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempyIntoNegCond4_G256_newbasis1);
    assign z6491_assgn6491 = dec_1_inp;
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> z2829_assgn2829);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z6497_assgn6497 = dec_1_inp;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & z2833_assgn2833);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z6503_assgn6503 = dec_11_inp;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ z2837_assgn2837);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempyIntoNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempyIntoNegCond5_G256_newbasis1);
    assign z6513_assgn6513 = dec_1_inp;
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> z2845_assgn2845);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z6519_assgn6519 = dec_1_inp;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & z2849_assgn2849);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z6525_assgn6525 = dec_158_inp;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ z2853_assgn2853);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempyIntoNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempyIntoNegCond6_G256_newbasis1);
    assign z6535_assgn6535 = dec_1_inp;
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> z2861_assgn2861);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z6541_assgn6541 = dec_1_inp;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & z2865_assgn2865);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z6547_assgn6547 = dec_45_inp;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ z2869_assgn2869);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempyIntoNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempyIntoNegCond7_G256_newbasis1);
    assign z6557_assgn6557 = dec_1_inp;
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> z2877_assgn2877);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z6563_assgn6563 = dec_1_inp;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & z2881_assgn2881);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z6569_assgn6569 = dec_88_inp;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ z2885_assgn2885);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempyIntoNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempyIntoNegCond8_G256_newbasis1);
    assign z6579_assgn6579 = dec_1_inp;
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> z2893_assgn2893);
    assign t7 = z_y8_G256_newbasis1;
    assign z6585_assgn6585 = dec_99_inp;

    always @(posedge clk) begin
        z3225_assgn32250 <= z3225_assgn3225;
        z3225_assgn32251 <= z3225_assgn32250;
        z3225_assgn32252 <= z3225_assgn32251;
        z3225_assgn32253 <= z3225_assgn32252;
        z3225_assgn32254 <= z3225_assgn32253;
        x8_G256_newbasis0 <= z3225_assgn32254;
        z3357_assgn33570 <= z3357_assgn3357;
        z3357_assgn33571 <= z3357_assgn33570;
        z3357_assgn33572 <= z3357_assgn33571;
        z3357_assgn33573 <= z3357_assgn33572;
        z3357_assgn33574 <= z3357_assgn33573;
        z_x8_G256_newbasis0 <= z3357_assgn33574;
        axorb_0_G4_mul0_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul0_G16_mul0_G256_inv0;
        b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= b1_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0;
        r10_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= r10_hpc10_G4_mul0_G16_mul0_G256_inv0;
        axorb_1_G4_mul0_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul0_G16_mul0_G256_inv0;
        b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= b0_preshared_hpc10_G4_mul0_G16_mul0_G256_inv0;
        i1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= i1_hpc10_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc10_G4_mul0_G16_mul0_G256_inv0;
        i2_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= i2_hpc10_G4_mul0_G16_mul0_G256_inv0;
        p4_hpc10_G4_mul0_G16_mul0_G256_inv0_reg <= p4_hpc10_G4_mul0_G16_mul0_G256_inv0;
        a0_G4_mul0_G16_mul0_G256_inv0_reg <= a0_G4_mul0_G16_mul0_G256_inv0;
        b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= b1_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0;
        r10_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= r10_hpc11_G4_mul0_G16_mul0_G256_inv0;
        a1_G4_mul0_G16_mul0_G256_inv0_reg <= a1_G4_mul0_G16_mul0_G256_inv0;
        b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= b0_preshared_hpc11_G4_mul0_G16_mul0_G256_inv0;
        i1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= i1_hpc11_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc11_G4_mul0_G16_mul0_G256_inv0;
        i2_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= i2_hpc11_G4_mul0_G16_mul0_G256_inv0;
        p4_hpc11_G4_mul0_G16_mul0_G256_inv0_reg <= p4_hpc11_G4_mul0_G16_mul0_G256_inv0;
        b0_G4_mul0_G16_mul0_G256_inv0_reg <= b0_G4_mul0_G16_mul0_G256_inv0;
        b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= b1_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0;
        r10_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= r10_hpc12_G4_mul0_G16_mul0_G256_inv0;
        b1_G4_mul0_G16_mul0_G256_inv0_reg <= b1_G4_mul0_G16_mul0_G256_inv0;
        b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= b0_preshared_hpc12_G4_mul0_G16_mul0_G256_inv0;
        i1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= i1_hpc12_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc12_G4_mul0_G16_mul0_G256_inv0;
        i2_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= i2_hpc12_G4_mul0_G16_mul0_G256_inv0;
        p4_hpc12_G4_mul0_G16_mul0_G256_inv0_reg <= p4_hpc12_G4_mul0_G16_mul0_G256_inv0;
        z3661_assgn36610 <= z3661_assgn3661;
        z761_assgn761 <= z3661_assgn36610;
        z3665_assgn36650 <= z3665_assgn3665;
        z763_assgn763 <= z3665_assgn36650;
        z3673_assgn36730 <= z3673_assgn3673;
        z769_assgn769 <= z3673_assgn36730;
        z3677_assgn36770 <= z3677_assgn3677;
        z771_assgn771 <= z3677_assgn36770;
        z3681_assgn36810 <= z3681_assgn3681;
        z773_assgn773 <= z3681_assgn36810;
        z3685_assgn36850 <= z3685_assgn3685;
        z775_assgn775 <= z3685_assgn36850;
        z3689_assgn36890 <= z3689_assgn3689;
        z777_assgn777 <= z3689_assgn36890;
        z3693_assgn36930 <= z3693_assgn3693;
        z779_assgn779 <= z3693_assgn36930;
        z3705_assgn37050 <= z3705_assgn3705;
        z789_assgn789 <= z3705_assgn37050;
        z3709_assgn37090 <= z3709_assgn3709;
        z791_assgn791 <= z3709_assgn37090;
        axorb_0_G4_mul1_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul1_G16_mul0_G256_inv0;
        b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= b1_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0;
        r10_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= r10_hpc10_G4_mul1_G16_mul0_G256_inv0;
        axorb_1_G4_mul1_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul1_G16_mul0_G256_inv0;
        b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= b0_preshared_hpc10_G4_mul1_G16_mul0_G256_inv0;
        i1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= i1_hpc10_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc10_G4_mul1_G16_mul0_G256_inv0;
        i2_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= i2_hpc10_G4_mul1_G16_mul0_G256_inv0;
        p4_hpc10_G4_mul1_G16_mul0_G256_inv0_reg <= p4_hpc10_G4_mul1_G16_mul0_G256_inv0;
        a0_G4_mul1_G16_mul0_G256_inv0_reg <= a0_G4_mul1_G16_mul0_G256_inv0;
        b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= b1_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0;
        r10_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= r10_hpc11_G4_mul1_G16_mul0_G256_inv0;
        a1_G4_mul1_G16_mul0_G256_inv0_reg <= a1_G4_mul1_G16_mul0_G256_inv0;
        b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= b0_preshared_hpc11_G4_mul1_G16_mul0_G256_inv0;
        i1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= i1_hpc11_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc11_G4_mul1_G16_mul0_G256_inv0;
        i2_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= i2_hpc11_G4_mul1_G16_mul0_G256_inv0;
        p4_hpc11_G4_mul1_G16_mul0_G256_inv0_reg <= p4_hpc11_G4_mul1_G16_mul0_G256_inv0;
        b0_G4_mul1_G16_mul0_G256_inv0_reg <= b0_G4_mul1_G16_mul0_G256_inv0;
        b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= b1_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0;
        r10_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= r10_hpc12_G4_mul1_G16_mul0_G256_inv0;
        b1_G4_mul1_G16_mul0_G256_inv0_reg <= b1_G4_mul1_G16_mul0_G256_inv0;
        b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= b0_preshared_hpc12_G4_mul1_G16_mul0_G256_inv0;
        i1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= i1_hpc12_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc12_G4_mul1_G16_mul0_G256_inv0;
        i2_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= i2_hpc12_G4_mul1_G16_mul0_G256_inv0;
        p4_hpc12_G4_mul1_G16_mul0_G256_inv0_reg <= p4_hpc12_G4_mul1_G16_mul0_G256_inv0;
        z3841_assgn38410 <= z3841_assgn3841;
        z921_assgn921 <= z3841_assgn38410;
        z3845_assgn38450 <= z3845_assgn3845;
        z923_assgn923 <= z3845_assgn38450;
        axorb_0_G4_mul2_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul2_G16_mul0_G256_inv0;
        b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= b1_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0;
        r10_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= r10_hpc10_G4_mul2_G16_mul0_G256_inv0;
        axorb_1_G4_mul2_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul2_G16_mul0_G256_inv0;
        b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= b0_preshared_hpc10_G4_mul2_G16_mul0_G256_inv0;
        i1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= i1_hpc10_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc10_G4_mul2_G16_mul0_G256_inv0;
        i2_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= i2_hpc10_G4_mul2_G16_mul0_G256_inv0;
        p4_hpc10_G4_mul2_G16_mul0_G256_inv0_reg <= p4_hpc10_G4_mul2_G16_mul0_G256_inv0;
        a0_G4_mul2_G16_mul0_G256_inv0_reg <= a0_G4_mul2_G16_mul0_G256_inv0;
        b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= b1_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0;
        r10_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= r10_hpc11_G4_mul2_G16_mul0_G256_inv0;
        a1_G4_mul2_G16_mul0_G256_inv0_reg <= a1_G4_mul2_G16_mul0_G256_inv0;
        b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= b0_preshared_hpc11_G4_mul2_G16_mul0_G256_inv0;
        i1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= i1_hpc11_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc11_G4_mul2_G16_mul0_G256_inv0;
        i2_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= i2_hpc11_G4_mul2_G16_mul0_G256_inv0;
        p4_hpc11_G4_mul2_G16_mul0_G256_inv0_reg <= p4_hpc11_G4_mul2_G16_mul0_G256_inv0;
        b0_G4_mul2_G16_mul0_G256_inv0_reg <= b0_G4_mul2_G16_mul0_G256_inv0;
        b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= b1_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0;
        r10_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= r10_hpc12_G4_mul2_G16_mul0_G256_inv0;
        b1_G4_mul2_G16_mul0_G256_inv0_reg <= b1_G4_mul2_G16_mul0_G256_inv0;
        b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= b0_preshared_hpc12_G4_mul2_G16_mul0_G256_inv0;
        i1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= i1_hpc12_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc12_G4_mul2_G16_mul0_G256_inv0;
        i2_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= i2_hpc12_G4_mul2_G16_mul0_G256_inv0;
        p4_hpc12_G4_mul2_G16_mul0_G256_inv0_reg <= p4_hpc12_G4_mul2_G16_mul0_G256_inv0;
        z3981_assgn39810 <= z3981_assgn3981;
        z1057_assgn1057 <= z3981_assgn39810;
        z3985_assgn39850 <= z3985_assgn3985;
        z1059_assgn1059 <= z3985_assgn39850;
        z3997_assgn39970 <= z3997_assgn3997;
        z1069_assgn1069 <= z3997_assgn39970;
        z4001_assgn40010 <= z4001_assgn4001;
        z1071_assgn1071 <= z4001_assgn40010;
        z4009_assgn40090 <= z4009_assgn4009;
        z1078_assgn1078 <= z4009_assgn40090;
        z4013_assgn40130 <= z4013_assgn4013;
        z1080_assgn1080 <= z4013_assgn40130;
        z4053_assgn40530 <= z4053_assgn4053;
        z1117_assgn1117 <= z4053_assgn40530;
        z4057_assgn40570 <= z4057_assgn4057;
        z1119_assgn1119 <= z4057_assgn40570;
        z4061_assgn40610 <= z4061_assgn4061;
        z1121_assgn1121 <= z4061_assgn40610;
        z4065_assgn40650 <= z4065_assgn4065;
        z1123_assgn1123 <= z4065_assgn40650;
        z4069_assgn40690 <= z4069_assgn4069;
        z1125_assgn1125 <= z4069_assgn40690;
        z4073_assgn40730 <= z4073_assgn4073;
        z1127_assgn1127 <= z4073_assgn40730;
        z4081_assgn40810 <= z4081_assgn4081;
        z1133_assgn1133 <= z4081_assgn40810;
        z4085_assgn40850 <= z4085_assgn4085;
        z1135_assgn1135 <= z4085_assgn40850;
        z4089_assgn40890 <= z4089_assgn4089;
        z1137_assgn1137 <= z4089_assgn40890;
        z4093_assgn40930 <= z4093_assgn4093;
        z1139_assgn1139 <= z4093_assgn40930;
        z4097_assgn40970 <= z4097_assgn4097;
        z1141_assgn1141 <= z4097_assgn40970;
        z4101_assgn41010 <= z4101_assgn4101;
        z1143_assgn1143 <= z4101_assgn41010;
        z4105_assgn41050 <= z4105_assgn4105;
        z1145_assgn1145 <= z4105_assgn41050;
        z4109_assgn41090 <= z4109_assgn4109;
        z1147_assgn1147 <= z4109_assgn41090;
        z4117_assgn41170 <= z4117_assgn4117;
        z1153_assgn1153 <= z4117_assgn41170;
        z4121_assgn41210 <= z4121_assgn4121;
        z1155_assgn1155 <= z4121_assgn41210;
        z4125_assgn41250 <= z4125_assgn4125;
        z1157_assgn1157 <= z4125_assgn41250;
        z4129_assgn41290 <= z4129_assgn4129;
        z1159_assgn1159 <= z4129_assgn41290;
        z4133_assgn41330 <= z4133_assgn4133;
        z1161_assgn1161 <= z4133_assgn41330;
        z4137_assgn41370 <= z4137_assgn4137;
        z1163_assgn1163 <= z4137_assgn41370;
        z4149_assgn41490 <= z4149_assgn4149;
        z1173_assgn1173 <= z4149_assgn41490;
        z4153_assgn41530 <= z4153_assgn4153;
        z1175_assgn1175 <= z4153_assgn41530;
        z4173_assgn41730 <= z4173_assgn4173;
        z1193_assgn1193 <= z4173_assgn41730;
        z4177_assgn41770 <= z4177_assgn4177;
        z1195_assgn1195 <= z4177_assgn41770;
        z4181_assgn41810 <= z4181_assgn4181;
        z1197_assgn1197 <= z4181_assgn41810;
        z4185_assgn41850 <= z4185_assgn4185;
        z1199_assgn1199 <= z4185_assgn41850;
        z4189_assgn41890 <= z4189_assgn4189;
        z1201_assgn1201 <= z4189_assgn41890;
        z4193_assgn41930 <= z4193_assgn4193;
        z1203_assgn1203 <= z4193_assgn41930;
        z4197_assgn41970 <= z4197_assgn4197;
        z1205_assgn1205 <= z4197_assgn41970;
        z4201_assgn42010 <= z4201_assgn4201;
        z1207_assgn1207 <= z4201_assgn42010;
        z4205_assgn42050 <= z4205_assgn4205;
        z1209_assgn1209 <= z4205_assgn42050;
        z4209_assgn42090 <= z4209_assgn4209;
        z1211_assgn1211 <= z4209_assgn42090;
        z4213_assgn42130 <= z4213_assgn4213;
        z1213_assgn1213 <= z4213_assgn42130;
        z4217_assgn42170 <= z4217_assgn4217;
        z1215_assgn1215 <= z4217_assgn42170;
        z4233_assgn42330 <= z4233_assgn4233;
        z1229_assgn1229 <= z4233_assgn42330;
        z4237_assgn42370 <= z4237_assgn4237;
        z1231_assgn1231 <= z4237_assgn42370;
        axorb_0_G4_mul3_G16_inv0_G256_inv0_reg <= axorb_0_G4_mul3_G16_inv0_G256_inv0;
        b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= b1_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0;
        z4243_assgn42430 <= z4243_assgn4243;
        z4243_assgn42431 <= z4243_assgn42430;
        z1235_assgn1235 <= z4243_assgn42431;
        axorb_1_G4_mul3_G16_inv0_G256_inv0_reg <= axorb_1_G4_mul3_G16_inv0_G256_inv0;
        b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= b0_preshared_hpc10_G4_mul3_G16_inv0_G256_inv0;
        z4249_assgn42490 <= z4249_assgn4249;
        z4249_assgn42491 <= z4249_assgn42490;
        z1239_assgn1239 <= z4249_assgn42491;
        i1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= i1_hpc10_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc10_G4_mul3_G16_inv0_G256_inv0;
        i2_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= i2_hpc10_G4_mul3_G16_inv0_G256_inv0;
        p4_hpc10_G4_mul3_G16_inv0_G256_inv0_reg <= p4_hpc10_G4_mul3_G16_inv0_G256_inv0;
        z4265_assgn42650 <= z4265_assgn4265;
        z1253_assgn1253 <= z4265_assgn42650;
        z4269_assgn42690 <= z4269_assgn4269;
        z1255_assgn1255 <= z4269_assgn42690;
        a0_G4_mul3_G16_inv0_G256_inv0_reg <= a0_G4_mul3_G16_inv0_G256_inv0;
        b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= b1_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0;
        z4275_assgn42750 <= z4275_assgn4275;
        z4275_assgn42751 <= z4275_assgn42750;
        z1259_assgn1259 <= z4275_assgn42751;
        a1_G4_mul3_G16_inv0_G256_inv0_reg <= a1_G4_mul3_G16_inv0_G256_inv0;
        b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= b0_preshared_hpc11_G4_mul3_G16_inv0_G256_inv0;
        z4281_assgn42810 <= z4281_assgn4281;
        z4281_assgn42811 <= z4281_assgn42810;
        z1263_assgn1263 <= z4281_assgn42811;
        i1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= i1_hpc11_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc11_G4_mul3_G16_inv0_G256_inv0;
        i2_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= i2_hpc11_G4_mul3_G16_inv0_G256_inv0;
        p4_hpc11_G4_mul3_G16_inv0_G256_inv0_reg <= p4_hpc11_G4_mul3_G16_inv0_G256_inv0;
        z4301_assgn43010 <= z4301_assgn4301;
        z1281_assgn1281 <= z4301_assgn43010;
        z4305_assgn43050 <= z4305_assgn4305;
        z1283_assgn1283 <= z4305_assgn43050;
        b0_G4_mul3_G16_inv0_G256_inv0_reg <= b0_G4_mul3_G16_inv0_G256_inv0;
        b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= b1_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0;
        z4311_assgn43110 <= z4311_assgn4311;
        z4311_assgn43111 <= z4311_assgn43110;
        z1287_assgn1287 <= z4311_assgn43111;
        b1_G4_mul3_G16_inv0_G256_inv0_reg <= b1_G4_mul3_G16_inv0_G256_inv0;
        b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= b0_preshared_hpc12_G4_mul3_G16_inv0_G256_inv0;
        z4317_assgn43170 <= z4317_assgn4317;
        z4317_assgn43171 <= z4317_assgn43170;
        z1291_assgn1291 <= z4317_assgn43171;
        i1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= i1_hpc12_G4_mul3_G16_inv0_G256_inv0;
        p1_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc12_G4_mul3_G16_inv0_G256_inv0;
        i2_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= i2_hpc12_G4_mul3_G16_inv0_G256_inv0;
        p4_hpc12_G4_mul3_G16_inv0_G256_inv0_reg <= p4_hpc12_G4_mul3_G16_inv0_G256_inv0;
        z4333_assgn43330 <= z4333_assgn4333;
        z4333_assgn43331 <= z4333_assgn43330;
        z4333_assgn43332 <= z4333_assgn43331;
        z1305_assgn1305 <= z4333_assgn43332;
        z4337_assgn43370 <= z4337_assgn4337;
        z4337_assgn43371 <= z4337_assgn43370;
        z4337_assgn43372 <= z4337_assgn43371;
        z1307_assgn1307 <= z4337_assgn43372;
        z4345_assgn43450 <= z4345_assgn4345;
        z1314_assgn1314 <= z4345_assgn43450;
        z4349_assgn43490 <= z4349_assgn4349;
        z1316_assgn1316 <= z4349_assgn43490;
        z4353_assgn43530 <= z4353_assgn4353;
        z4353_assgn43531 <= z4353_assgn43530;
        z4353_assgn43532 <= z4353_assgn43531;
        z1317_assgn1317 <= z4353_assgn43532;
        z4357_assgn43570 <= z4357_assgn4357;
        z4357_assgn43571 <= z4357_assgn43570;
        z4357_assgn43572 <= z4357_assgn43571;
        z1319_assgn1319 <= z4357_assgn43572;
        z4361_assgn43610 <= z4361_assgn4361;
        z4361_assgn43611 <= z4361_assgn43610;
        z4361_assgn43612 <= z4361_assgn43611;
        z1321_assgn1321 <= z4361_assgn43612;
        z4365_assgn43650 <= z4365_assgn4365;
        z4365_assgn43651 <= z4365_assgn43650;
        z4365_assgn43652 <= z4365_assgn43651;
        z1323_assgn1323 <= z4365_assgn43652;
        z4369_assgn43690 <= z4369_assgn4369;
        z4369_assgn43691 <= z4369_assgn43690;
        z4369_assgn43692 <= z4369_assgn43691;
        z1325_assgn1325 <= z4369_assgn43692;
        z4373_assgn43730 <= z4373_assgn4373;
        z4373_assgn43731 <= z4373_assgn43730;
        z4373_assgn43732 <= z4373_assgn43731;
        z1327_assgn1327 <= z4373_assgn43732;
        z4377_assgn43770 <= z4377_assgn4377;
        z4377_assgn43771 <= z4377_assgn43770;
        z4377_assgn43772 <= z4377_assgn43771;
        z1329_assgn1329 <= z4377_assgn43772;
        z4381_assgn43810 <= z4381_assgn4381;
        z4381_assgn43811 <= z4381_assgn43810;
        z4381_assgn43812 <= z4381_assgn43811;
        z1331_assgn1331 <= z4381_assgn43812;
        z4401_assgn44010 <= z4401_assgn4401;
        z4401_assgn44011 <= z4401_assgn44010;
        z4401_assgn44012 <= z4401_assgn44011;
        z1349_assgn1349 <= z4401_assgn44012;
        z4405_assgn44050 <= z4405_assgn4405;
        z4405_assgn44051 <= z4405_assgn44050;
        z4405_assgn44052 <= z4405_assgn44051;
        z1351_assgn1351 <= z4405_assgn44052;
        z4409_assgn44090 <= z4409_assgn4409;
        z4409_assgn44091 <= z4409_assgn44090;
        z4409_assgn44092 <= z4409_assgn44091;
        z1353_assgn1353 <= z4409_assgn44092;
        z4413_assgn44130 <= z4413_assgn4413;
        z4413_assgn44131 <= z4413_assgn44130;
        z4413_assgn44132 <= z4413_assgn44131;
        z1355_assgn1355 <= z4413_assgn44132;
        z4417_assgn44170 <= z4417_assgn4417;
        z4417_assgn44171 <= z4417_assgn44170;
        z4417_assgn44172 <= z4417_assgn44171;
        z1357_assgn1357 <= z4417_assgn44172;
        z4421_assgn44210 <= z4421_assgn4421;
        z4421_assgn44211 <= z4421_assgn44210;
        z4421_assgn44212 <= z4421_assgn44211;
        z1359_assgn1359 <= z4421_assgn44212;
        z4425_assgn44250 <= z4425_assgn4425;
        z1361_assgn1361 <= z4425_assgn44250;
        z4429_assgn44290 <= z4429_assgn4429;
        z1363_assgn1363 <= z4429_assgn44290;
        z4433_assgn44330 <= z4433_assgn4433;
        z1365_assgn1365 <= z4433_assgn44330;
        z4437_assgn44370 <= z4437_assgn4437;
        z1367_assgn1367 <= z4437_assgn44370;
        z4441_assgn44410 <= z4441_assgn4441;
        z1369_assgn1369 <= z4441_assgn44410;
        z4445_assgn44450 <= z4445_assgn4445;
        z1371_assgn1371 <= z4445_assgn44450;
        z4461_assgn44610 <= z4461_assgn4461;
        z1385_assgn1385 <= z4461_assgn44610;
        z4465_assgn44650 <= z4465_assgn4465;
        z1387_assgn1387 <= z4465_assgn44650;
        z4469_assgn44690 <= z4469_assgn4469;
        z1389_assgn1389 <= z4469_assgn44690;
        z4473_assgn44730 <= z4473_assgn4473;
        z4473_assgn44731 <= z4473_assgn44730;
        z4473_assgn44732 <= z4473_assgn44731;
        z1391_assgn1391 <= z4473_assgn44732;
        z4477_assgn44770 <= z4477_assgn4477;
        z1393_assgn1393 <= z4477_assgn44770;
        z4481_assgn44810 <= z4481_assgn4481;
        z4481_assgn44811 <= z4481_assgn44810;
        z4481_assgn44812 <= z4481_assgn44811;
        z1395_assgn1395 <= z4481_assgn44812;
        z4485_assgn44850 <= z4485_assgn4485;
        z1397_assgn1397 <= z4485_assgn44850;
        z4489_assgn44890 <= z4489_assgn4489;
        z1399_assgn1399 <= z4489_assgn44890;
        i1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg <= i1_hpc10_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc10_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc10_G4_mul4_G16_inv0_G256_inv0;
        i2_hpc10_G4_mul4_G16_inv0_G256_inv0_reg <= i2_hpc10_G4_mul4_G16_inv0_G256_inv0;
        p4_hpc10_G4_mul4_G16_inv0_G256_inv0_reg <= p4_hpc10_G4_mul4_G16_inv0_G256_inv0;
        z4501_assgn45010 <= z4501_assgn4501;
        z1409_assgn1409 <= z4501_assgn45010;
        z4505_assgn45050 <= z4505_assgn4505;
        z1411_assgn1411 <= z4505_assgn45050;
        z4509_assgn45090 <= z4509_assgn4509;
        z1413_assgn1413 <= z4509_assgn45090;
        z4513_assgn45130 <= z4513_assgn4513;
        z4513_assgn45131 <= z4513_assgn45130;
        z4513_assgn45132 <= z4513_assgn45131;
        z1415_assgn1415 <= z4513_assgn45132;
        z4517_assgn45170 <= z4517_assgn4517;
        z1417_assgn1417 <= z4517_assgn45170;
        z4521_assgn45210 <= z4521_assgn4521;
        z4521_assgn45211 <= z4521_assgn45210;
        z4521_assgn45212 <= z4521_assgn45211;
        z1419_assgn1419 <= z4521_assgn45212;
        z4525_assgn45250 <= z4525_assgn4525;
        z1421_assgn1421 <= z4525_assgn45250;
        z4529_assgn45290 <= z4529_assgn4529;
        z1423_assgn1423 <= z4529_assgn45290;
        i1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg <= i1_hpc11_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc11_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc11_G4_mul4_G16_inv0_G256_inv0;
        i2_hpc11_G4_mul4_G16_inv0_G256_inv0_reg <= i2_hpc11_G4_mul4_G16_inv0_G256_inv0;
        p4_hpc11_G4_mul4_G16_inv0_G256_inv0_reg <= p4_hpc11_G4_mul4_G16_inv0_G256_inv0;
        z4545_assgn45450 <= z4545_assgn4545;
        z1437_assgn1437 <= z4545_assgn45450;
        z4549_assgn45490 <= z4549_assgn4549;
        z1439_assgn1439 <= z4549_assgn45490;
        z4553_assgn45530 <= z4553_assgn4553;
        z1441_assgn1441 <= z4553_assgn45530;
        z4557_assgn45570 <= z4557_assgn4557;
        z4557_assgn45571 <= z4557_assgn45570;
        z4557_assgn45572 <= z4557_assgn45571;
        z1443_assgn1443 <= z4557_assgn45572;
        z4561_assgn45610 <= z4561_assgn4561;
        z1445_assgn1445 <= z4561_assgn45610;
        z4565_assgn45650 <= z4565_assgn4565;
        z4565_assgn45651 <= z4565_assgn45650;
        z4565_assgn45652 <= z4565_assgn45651;
        z1447_assgn1447 <= z4565_assgn45652;
        z4569_assgn45690 <= z4569_assgn4569;
        z1449_assgn1449 <= z4569_assgn45690;
        z4573_assgn45730 <= z4573_assgn4573;
        z1451_assgn1451 <= z4573_assgn45730;
        i1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg <= i1_hpc12_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc12_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc12_G4_mul4_G16_inv0_G256_inv0;
        i2_hpc12_G4_mul4_G16_inv0_G256_inv0_reg <= i2_hpc12_G4_mul4_G16_inv0_G256_inv0;
        p4_hpc12_G4_mul4_G16_inv0_G256_inv0_reg <= p4_hpc12_G4_mul4_G16_inv0_G256_inv0;
        z4585_assgn45850 <= z4585_assgn4585;
        z4585_assgn45851 <= z4585_assgn45850;
        z4585_assgn45852 <= z4585_assgn45851;
        z4585_assgn45853 <= z4585_assgn45852;
        z1461_assgn1461 <= z4585_assgn45853;
        z4589_assgn45890 <= z4589_assgn4589;
        z4589_assgn45891 <= z4589_assgn45890;
        z4589_assgn45892 <= z4589_assgn45891;
        z4589_assgn45893 <= z4589_assgn45892;
        z1463_assgn1463 <= z4589_assgn45893;
        z4609_assgn46090 <= z4609_assgn4609;
        z4609_assgn46091 <= z4609_assgn46090;
        z4609_assgn46092 <= z4609_assgn46091;
        z1481_assgn1481 <= z4609_assgn46092;
        z4613_assgn46130 <= z4613_assgn4613;
        z4613_assgn46131 <= z4613_assgn46130;
        z4613_assgn46132 <= z4613_assgn46131;
        z1483_assgn1483 <= z4613_assgn46132;
        z4617_assgn46170 <= z4617_assgn4617;
        z4617_assgn46171 <= z4617_assgn46170;
        z4617_assgn46172 <= z4617_assgn46171;
        z1485_assgn1485 <= z4617_assgn46172;
        z4621_assgn46210 <= z4621_assgn4621;
        z4621_assgn46211 <= z4621_assgn46210;
        z4621_assgn46212 <= z4621_assgn46211;
        z1487_assgn1487 <= z4621_assgn46212;
        z4625_assgn46250 <= z4625_assgn4625;
        z4625_assgn46251 <= z4625_assgn46250;
        z4625_assgn46252 <= z4625_assgn46251;
        z1489_assgn1489 <= z4625_assgn46252;
        z4629_assgn46290 <= z4629_assgn4629;
        z4629_assgn46291 <= z4629_assgn46290;
        z4629_assgn46292 <= z4629_assgn46291;
        z1491_assgn1491 <= z4629_assgn46292;
        z4633_assgn46330 <= z4633_assgn4633;
        z1493_assgn1493 <= z4633_assgn46330;
        z4637_assgn46370 <= z4637_assgn4637;
        z1495_assgn1495 <= z4637_assgn46370;
        z4641_assgn46410 <= z4641_assgn4641;
        z1497_assgn1497 <= z4641_assgn46410;
        z4645_assgn46450 <= z4645_assgn4645;
        z1499_assgn1499 <= z4645_assgn46450;
        z4649_assgn46490 <= z4649_assgn4649;
        z1501_assgn1501 <= z4649_assgn46490;
        z4653_assgn46530 <= z4653_assgn4653;
        z1503_assgn1503 <= z4653_assgn46530;
        z4669_assgn46690 <= z4669_assgn4669;
        z1517_assgn1517 <= z4669_assgn46690;
        z4673_assgn46730 <= z4673_assgn4673;
        z1519_assgn1519 <= z4673_assgn46730;
        z4677_assgn46770 <= z4677_assgn4677;
        z1521_assgn1521 <= z4677_assgn46770;
        z4681_assgn46810 <= z4681_assgn4681;
        z4681_assgn46811 <= z4681_assgn46810;
        z4681_assgn46812 <= z4681_assgn46811;
        z1523_assgn1523 <= z4681_assgn46812;
        z4685_assgn46850 <= z4685_assgn4685;
        z1525_assgn1525 <= z4685_assgn46850;
        z4689_assgn46890 <= z4689_assgn4689;
        z4689_assgn46891 <= z4689_assgn46890;
        z4689_assgn46892 <= z4689_assgn46891;
        z1527_assgn1527 <= z4689_assgn46892;
        z4693_assgn46930 <= z4693_assgn4693;
        z1529_assgn1529 <= z4693_assgn46930;
        z4697_assgn46970 <= z4697_assgn4697;
        z1531_assgn1531 <= z4697_assgn46970;
        i1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg <= i1_hpc10_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc10_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc10_G4_mul5_G16_inv0_G256_inv0;
        i2_hpc10_G4_mul5_G16_inv0_G256_inv0_reg <= i2_hpc10_G4_mul5_G16_inv0_G256_inv0;
        p4_hpc10_G4_mul5_G16_inv0_G256_inv0_reg <= p4_hpc10_G4_mul5_G16_inv0_G256_inv0;
        z4709_assgn47090 <= z4709_assgn4709;
        z1541_assgn1541 <= z4709_assgn47090;
        z4713_assgn47130 <= z4713_assgn4713;
        z1543_assgn1543 <= z4713_assgn47130;
        z4717_assgn47170 <= z4717_assgn4717;
        z1545_assgn1545 <= z4717_assgn47170;
        z4721_assgn47210 <= z4721_assgn4721;
        z4721_assgn47211 <= z4721_assgn47210;
        z4721_assgn47212 <= z4721_assgn47211;
        z1547_assgn1547 <= z4721_assgn47212;
        z4725_assgn47250 <= z4725_assgn4725;
        z1549_assgn1549 <= z4725_assgn47250;
        z4729_assgn47290 <= z4729_assgn4729;
        z4729_assgn47291 <= z4729_assgn47290;
        z4729_assgn47292 <= z4729_assgn47291;
        z1551_assgn1551 <= z4729_assgn47292;
        z4733_assgn47330 <= z4733_assgn4733;
        z1553_assgn1553 <= z4733_assgn47330;
        z4737_assgn47370 <= z4737_assgn4737;
        z1555_assgn1555 <= z4737_assgn47370;
        i1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg <= i1_hpc11_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc11_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc11_G4_mul5_G16_inv0_G256_inv0;
        i2_hpc11_G4_mul5_G16_inv0_G256_inv0_reg <= i2_hpc11_G4_mul5_G16_inv0_G256_inv0;
        p4_hpc11_G4_mul5_G16_inv0_G256_inv0_reg <= p4_hpc11_G4_mul5_G16_inv0_G256_inv0;
        z4753_assgn47530 <= z4753_assgn4753;
        z1569_assgn1569 <= z4753_assgn47530;
        z4757_assgn47570 <= z4757_assgn4757;
        z1571_assgn1571 <= z4757_assgn47570;
        z4761_assgn47610 <= z4761_assgn4761;
        z1573_assgn1573 <= z4761_assgn47610;
        z4765_assgn47650 <= z4765_assgn4765;
        z4765_assgn47651 <= z4765_assgn47650;
        z4765_assgn47652 <= z4765_assgn47651;
        z1575_assgn1575 <= z4765_assgn47652;
        z4769_assgn47690 <= z4769_assgn4769;
        z1577_assgn1577 <= z4769_assgn47690;
        z4773_assgn47730 <= z4773_assgn4773;
        z4773_assgn47731 <= z4773_assgn47730;
        z4773_assgn47732 <= z4773_assgn47731;
        z1579_assgn1579 <= z4773_assgn47732;
        z4777_assgn47770 <= z4777_assgn4777;
        z1581_assgn1581 <= z4777_assgn47770;
        z4781_assgn47810 <= z4781_assgn4781;
        z1583_assgn1583 <= z4781_assgn47810;
        i1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg <= i1_hpc12_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc12_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc12_G4_mul5_G16_inv0_G256_inv0;
        i2_hpc12_G4_mul5_G16_inv0_G256_inv0_reg <= i2_hpc12_G4_mul5_G16_inv0_G256_inv0;
        p4_hpc12_G4_mul5_G16_inv0_G256_inv0_reg <= p4_hpc12_G4_mul5_G16_inv0_G256_inv0;
        z4793_assgn47930 <= z4793_assgn4793;
        z4793_assgn47931 <= z4793_assgn47930;
        z4793_assgn47932 <= z4793_assgn47931;
        z4793_assgn47933 <= z4793_assgn47932;
        z1593_assgn1593 <= z4793_assgn47933;
        z4797_assgn47970 <= z4797_assgn4797;
        z4797_assgn47971 <= z4797_assgn47970;
        z4797_assgn47972 <= z4797_assgn47971;
        z4797_assgn47973 <= z4797_assgn47972;
        z1595_assgn1595 <= z4797_assgn47973;
        z4805_assgn48050 <= z4805_assgn4805;
        z4805_assgn48051 <= z4805_assgn48050;
        z4805_assgn48052 <= z4805_assgn48051;
        z4805_assgn48053 <= z4805_assgn48052;
        z1601_assgn1601 <= z4805_assgn48053;
        z4809_assgn48090 <= z4809_assgn4809;
        z4809_assgn48091 <= z4809_assgn48090;
        z4809_assgn48092 <= z4809_assgn48091;
        z4809_assgn48093 <= z4809_assgn48092;
        z1603_assgn1603 <= z4809_assgn48093;
        z4853_assgn48530 <= z4853_assgn4853;
        z4853_assgn48531 <= z4853_assgn48530;
        z4853_assgn48532 <= z4853_assgn48531;
        z4853_assgn48533 <= z4853_assgn48532;
        z1645_assgn1645 <= z4853_assgn48533;
        z4857_assgn48570 <= z4857_assgn4857;
        z4857_assgn48571 <= z4857_assgn48570;
        z4857_assgn48572 <= z4857_assgn48571;
        z4857_assgn48573 <= z4857_assgn48572;
        z1647_assgn1647 <= z4857_assgn48573;
        z4861_assgn48610 <= z4861_assgn4861;
        z4861_assgn48611 <= z4861_assgn48610;
        z4861_assgn48612 <= z4861_assgn48611;
        z4861_assgn48613 <= z4861_assgn48612;
        z1649_assgn1649 <= z4861_assgn48613;
        z4865_assgn48650 <= z4865_assgn4865;
        z4865_assgn48651 <= z4865_assgn48650;
        z4865_assgn48652 <= z4865_assgn48651;
        z4865_assgn48653 <= z4865_assgn48652;
        z1651_assgn1651 <= z4865_assgn48653;
        z4869_assgn48690 <= z4869_assgn4869;
        z4869_assgn48691 <= z4869_assgn48690;
        z4869_assgn48692 <= z4869_assgn48691;
        z4869_assgn48693 <= z4869_assgn48692;
        z1653_assgn1653 <= z4869_assgn48693;
        z4873_assgn48730 <= z4873_assgn4873;
        z4873_assgn48731 <= z4873_assgn48730;
        z4873_assgn48732 <= z4873_assgn48731;
        z4873_assgn48733 <= z4873_assgn48732;
        z1655_assgn1655 <= z4873_assgn48733;
        z4909_assgn49090 <= z4909_assgn4909;
        z4909_assgn49091 <= z4909_assgn49090;
        z4909_assgn49092 <= z4909_assgn49091;
        z4909_assgn49093 <= z4909_assgn49092;
        z1689_assgn1689 <= z4909_assgn49093;
        z4913_assgn49130 <= z4913_assgn4913;
        z4913_assgn49131 <= z4913_assgn49130;
        z4913_assgn49132 <= z4913_assgn49131;
        z4913_assgn49133 <= z4913_assgn49132;
        z1691_assgn1691 <= z4913_assgn49133;
        z4917_assgn49170 <= z4917_assgn4917;
        z4917_assgn49171 <= z4917_assgn49170;
        z4917_assgn49172 <= z4917_assgn49171;
        z4917_assgn49173 <= z4917_assgn49172;
        z1693_assgn1693 <= z4917_assgn49173;
        z4921_assgn49210 <= z4921_assgn4921;
        z4921_assgn49211 <= z4921_assgn49210;
        z4921_assgn49212 <= z4921_assgn49211;
        z4921_assgn49213 <= z4921_assgn49212;
        z1695_assgn1695 <= z4921_assgn49213;
        z4925_assgn49250 <= z4925_assgn4925;
        z4925_assgn49251 <= z4925_assgn49250;
        z4925_assgn49252 <= z4925_assgn49251;
        z4925_assgn49253 <= z4925_assgn49252;
        z1697_assgn1697 <= z4925_assgn49253;
        z4929_assgn49290 <= z4929_assgn4929;
        z4929_assgn49291 <= z4929_assgn49290;
        z4929_assgn49292 <= z4929_assgn49291;
        z4929_assgn49293 <= z4929_assgn49292;
        z1699_assgn1699 <= z4929_assgn49293;
        z4961_assgn49610 <= z4961_assgn4961;
        z4961_assgn49611 <= z4961_assgn49610;
        z4961_assgn49612 <= z4961_assgn49611;
        z4961_assgn49613 <= z4961_assgn49612;
        z1729_assgn1729 <= z4961_assgn49613;
        z4965_assgn49650 <= z4965_assgn4965;
        z4965_assgn49651 <= z4965_assgn49650;
        z4965_assgn49652 <= z4965_assgn49651;
        z4965_assgn49653 <= z4965_assgn49652;
        z1731_assgn1731 <= z4965_assgn49653;
        z4969_assgn49690 <= z4969_assgn4969;
        z4969_assgn49691 <= z4969_assgn49690;
        z4969_assgn49692 <= z4969_assgn49691;
        z4969_assgn49693 <= z4969_assgn49692;
        z1733_assgn1733 <= z4969_assgn49693;
        z4973_assgn49730 <= z4973_assgn4973;
        z4973_assgn49731 <= z4973_assgn49730;
        z4973_assgn49732 <= z4973_assgn49731;
        z4973_assgn49733 <= z4973_assgn49732;
        z1735_assgn1735 <= z4973_assgn49733;
        z4977_assgn49770 <= z4977_assgn4977;
        z4977_assgn49771 <= z4977_assgn49770;
        z4977_assgn49772 <= z4977_assgn49771;
        z4977_assgn49773 <= z4977_assgn49772;
        z1737_assgn1737 <= z4977_assgn49773;
        z4981_assgn49810 <= z4981_assgn4981;
        z4981_assgn49811 <= z4981_assgn49810;
        z4981_assgn49812 <= z4981_assgn49811;
        z4981_assgn49813 <= z4981_assgn49812;
        z1739_assgn1739 <= z4981_assgn49813;
        i1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg <= i1_hpc10_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc10_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc10_G4_mul0_G16_mul1_G256_inv0;
        i2_hpc10_G4_mul0_G16_mul1_G256_inv0_reg <= i2_hpc10_G4_mul0_G16_mul1_G256_inv0;
        p4_hpc10_G4_mul0_G16_mul1_G256_inv0_reg <= p4_hpc10_G4_mul0_G16_mul1_G256_inv0;
        z4997_assgn49970 <= z4997_assgn4997;
        z4997_assgn49971 <= z4997_assgn49970;
        z4997_assgn49972 <= z4997_assgn49971;
        z4997_assgn49973 <= z4997_assgn49972;
        z1753_assgn1753 <= z4997_assgn49973;
        z5001_assgn50010 <= z5001_assgn5001;
        z5001_assgn50011 <= z5001_assgn50010;
        z5001_assgn50012 <= z5001_assgn50011;
        z5001_assgn50013 <= z5001_assgn50012;
        z1755_assgn1755 <= z5001_assgn50013;
        z5005_assgn50050 <= z5005_assgn5005;
        z5005_assgn50051 <= z5005_assgn50050;
        z5005_assgn50052 <= z5005_assgn50051;
        z5005_assgn50053 <= z5005_assgn50052;
        z1757_assgn1757 <= z5005_assgn50053;
        z5009_assgn50090 <= z5009_assgn5009;
        z5009_assgn50091 <= z5009_assgn50090;
        z5009_assgn50092 <= z5009_assgn50091;
        z5009_assgn50093 <= z5009_assgn50092;
        z1759_assgn1759 <= z5009_assgn50093;
        z5013_assgn50130 <= z5013_assgn5013;
        z5013_assgn50131 <= z5013_assgn50130;
        z5013_assgn50132 <= z5013_assgn50131;
        z5013_assgn50133 <= z5013_assgn50132;
        z1761_assgn1761 <= z5013_assgn50133;
        z5017_assgn50170 <= z5017_assgn5017;
        z5017_assgn50171 <= z5017_assgn50170;
        z5017_assgn50172 <= z5017_assgn50171;
        z5017_assgn50173 <= z5017_assgn50172;
        z1763_assgn1763 <= z5017_assgn50173;
        i1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg <= i1_hpc11_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc11_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc11_G4_mul0_G16_mul1_G256_inv0;
        i2_hpc11_G4_mul0_G16_mul1_G256_inv0_reg <= i2_hpc11_G4_mul0_G16_mul1_G256_inv0;
        p4_hpc11_G4_mul0_G16_mul1_G256_inv0_reg <= p4_hpc11_G4_mul0_G16_mul1_G256_inv0;
        z5037_assgn50370 <= z5037_assgn5037;
        z5037_assgn50371 <= z5037_assgn50370;
        z5037_assgn50372 <= z5037_assgn50371;
        z5037_assgn50373 <= z5037_assgn50372;
        z1781_assgn1781 <= z5037_assgn50373;
        z5041_assgn50410 <= z5041_assgn5041;
        z5041_assgn50411 <= z5041_assgn50410;
        z5041_assgn50412 <= z5041_assgn50411;
        z5041_assgn50413 <= z5041_assgn50412;
        z1783_assgn1783 <= z5041_assgn50413;
        z5045_assgn50450 <= z5045_assgn5045;
        z5045_assgn50451 <= z5045_assgn50450;
        z5045_assgn50452 <= z5045_assgn50451;
        z5045_assgn50453 <= z5045_assgn50452;
        z1785_assgn1785 <= z5045_assgn50453;
        z5049_assgn50490 <= z5049_assgn5049;
        z5049_assgn50491 <= z5049_assgn50490;
        z5049_assgn50492 <= z5049_assgn50491;
        z5049_assgn50493 <= z5049_assgn50492;
        z1787_assgn1787 <= z5049_assgn50493;
        z5053_assgn50530 <= z5053_assgn5053;
        z5053_assgn50531 <= z5053_assgn50530;
        z5053_assgn50532 <= z5053_assgn50531;
        z5053_assgn50533 <= z5053_assgn50532;
        z1789_assgn1789 <= z5053_assgn50533;
        z5057_assgn50570 <= z5057_assgn5057;
        z5057_assgn50571 <= z5057_assgn50570;
        z5057_assgn50572 <= z5057_assgn50571;
        z5057_assgn50573 <= z5057_assgn50572;
        z1791_assgn1791 <= z5057_assgn50573;
        i1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg <= i1_hpc12_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc12_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc12_G4_mul0_G16_mul1_G256_inv0;
        i2_hpc12_G4_mul0_G16_mul1_G256_inv0_reg <= i2_hpc12_G4_mul0_G16_mul1_G256_inv0;
        p4_hpc12_G4_mul0_G16_mul1_G256_inv0_reg <= p4_hpc12_G4_mul0_G16_mul1_G256_inv0;
        z5069_assgn50690 <= z5069_assgn5069;
        z5069_assgn50691 <= z5069_assgn50690;
        z5069_assgn50692 <= z5069_assgn50691;
        z5069_assgn50693 <= z5069_assgn50692;
        z5069_assgn50694 <= z5069_assgn50693;
        z1801_assgn1801 <= z5069_assgn50694;
        z5073_assgn50730 <= z5073_assgn5073;
        z5073_assgn50731 <= z5073_assgn50730;
        z5073_assgn50732 <= z5073_assgn50731;
        z5073_assgn50733 <= z5073_assgn50732;
        z5073_assgn50734 <= z5073_assgn50733;
        z1803_assgn1803 <= z5073_assgn50734;
        z5081_assgn50810 <= z5081_assgn5081;
        z5081_assgn50811 <= z5081_assgn50810;
        z5081_assgn50812 <= z5081_assgn50811;
        z5081_assgn50813 <= z5081_assgn50812;
        z5081_assgn50814 <= z5081_assgn50813;
        z1809_assgn1809 <= z5081_assgn50814;
        z5085_assgn50850 <= z5085_assgn5085;
        z5085_assgn50851 <= z5085_assgn50850;
        z5085_assgn50852 <= z5085_assgn50851;
        z5085_assgn50853 <= z5085_assgn50852;
        z5085_assgn50854 <= z5085_assgn50853;
        z1811_assgn1811 <= z5085_assgn50854;
        z5089_assgn50890 <= z5089_assgn5089;
        z5089_assgn50891 <= z5089_assgn50890;
        z5089_assgn50892 <= z5089_assgn50891;
        z5089_assgn50893 <= z5089_assgn50892;
        z5089_assgn50894 <= z5089_assgn50893;
        z1813_assgn1813 <= z5089_assgn50894;
        z5093_assgn50930 <= z5093_assgn5093;
        z5093_assgn50931 <= z5093_assgn50930;
        z5093_assgn50932 <= z5093_assgn50931;
        z5093_assgn50933 <= z5093_assgn50932;
        z5093_assgn50934 <= z5093_assgn50933;
        z1815_assgn1815 <= z5093_assgn50934;
        z5097_assgn50970 <= z5097_assgn5097;
        z5097_assgn50971 <= z5097_assgn50970;
        z5097_assgn50972 <= z5097_assgn50971;
        z5097_assgn50973 <= z5097_assgn50972;
        z5097_assgn50974 <= z5097_assgn50973;
        z1817_assgn1817 <= z5097_assgn50974;
        z5101_assgn51010 <= z5101_assgn5101;
        z5101_assgn51011 <= z5101_assgn51010;
        z5101_assgn51012 <= z5101_assgn51011;
        z5101_assgn51013 <= z5101_assgn51012;
        z5101_assgn51014 <= z5101_assgn51013;
        z1819_assgn1819 <= z5101_assgn51014;
        z5113_assgn51130 <= z5113_assgn5113;
        z5113_assgn51131 <= z5113_assgn51130;
        z5113_assgn51132 <= z5113_assgn51131;
        z5113_assgn51133 <= z5113_assgn51132;
        z5113_assgn51134 <= z5113_assgn51133;
        z1829_assgn1829 <= z5113_assgn51134;
        z5117_assgn51170 <= z5117_assgn5117;
        z5117_assgn51171 <= z5117_assgn51170;
        z5117_assgn51172 <= z5117_assgn51171;
        z5117_assgn51173 <= z5117_assgn51172;
        z5117_assgn51174 <= z5117_assgn51173;
        z1831_assgn1831 <= z5117_assgn51174;
        z5137_assgn51370 <= z5137_assgn5137;
        z5137_assgn51371 <= z5137_assgn51370;
        z5137_assgn51372 <= z5137_assgn51371;
        z5137_assgn51373 <= z5137_assgn51372;
        z1849_assgn1849 <= z5137_assgn51373;
        z5141_assgn51410 <= z5141_assgn5141;
        z5141_assgn51411 <= z5141_assgn51410;
        z5141_assgn51412 <= z5141_assgn51411;
        z5141_assgn51413 <= z5141_assgn51412;
        z1851_assgn1851 <= z5141_assgn51413;
        z5145_assgn51450 <= z5145_assgn5145;
        z5145_assgn51451 <= z5145_assgn51450;
        z5145_assgn51452 <= z5145_assgn51451;
        z5145_assgn51453 <= z5145_assgn51452;
        z1853_assgn1853 <= z5145_assgn51453;
        z5149_assgn51490 <= z5149_assgn5149;
        z5149_assgn51491 <= z5149_assgn51490;
        z5149_assgn51492 <= z5149_assgn51491;
        z5149_assgn51493 <= z5149_assgn51492;
        z1855_assgn1855 <= z5149_assgn51493;
        z5153_assgn51530 <= z5153_assgn5153;
        z5153_assgn51531 <= z5153_assgn51530;
        z5153_assgn51532 <= z5153_assgn51531;
        z5153_assgn51533 <= z5153_assgn51532;
        z1857_assgn1857 <= z5153_assgn51533;
        z5157_assgn51570 <= z5157_assgn5157;
        z5157_assgn51571 <= z5157_assgn51570;
        z5157_assgn51572 <= z5157_assgn51571;
        z5157_assgn51573 <= z5157_assgn51572;
        z1859_assgn1859 <= z5157_assgn51573;
        z5189_assgn51890 <= z5189_assgn5189;
        z5189_assgn51891 <= z5189_assgn51890;
        z5189_assgn51892 <= z5189_assgn51891;
        z5189_assgn51893 <= z5189_assgn51892;
        z1889_assgn1889 <= z5189_assgn51893;
        z5193_assgn51930 <= z5193_assgn5193;
        z5193_assgn51931 <= z5193_assgn51930;
        z5193_assgn51932 <= z5193_assgn51931;
        z5193_assgn51933 <= z5193_assgn51932;
        z1891_assgn1891 <= z5193_assgn51933;
        z5197_assgn51970 <= z5197_assgn5197;
        z5197_assgn51971 <= z5197_assgn51970;
        z5197_assgn51972 <= z5197_assgn51971;
        z5197_assgn51973 <= z5197_assgn51972;
        z1893_assgn1893 <= z5197_assgn51973;
        z5201_assgn52010 <= z5201_assgn5201;
        z5201_assgn52011 <= z5201_assgn52010;
        z5201_assgn52012 <= z5201_assgn52011;
        z5201_assgn52013 <= z5201_assgn52012;
        z1895_assgn1895 <= z5201_assgn52013;
        z5205_assgn52050 <= z5205_assgn5205;
        z5205_assgn52051 <= z5205_assgn52050;
        z5205_assgn52052 <= z5205_assgn52051;
        z5205_assgn52053 <= z5205_assgn52052;
        z1897_assgn1897 <= z5205_assgn52053;
        z5209_assgn52090 <= z5209_assgn5209;
        z5209_assgn52091 <= z5209_assgn52090;
        z5209_assgn52092 <= z5209_assgn52091;
        z5209_assgn52093 <= z5209_assgn52092;
        z1899_assgn1899 <= z5209_assgn52093;
        i1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg <= i1_hpc10_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc10_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc10_G4_mul1_G16_mul1_G256_inv0;
        i2_hpc10_G4_mul1_G16_mul1_G256_inv0_reg <= i2_hpc10_G4_mul1_G16_mul1_G256_inv0;
        p4_hpc10_G4_mul1_G16_mul1_G256_inv0_reg <= p4_hpc10_G4_mul1_G16_mul1_G256_inv0;
        z5225_assgn52250 <= z5225_assgn5225;
        z5225_assgn52251 <= z5225_assgn52250;
        z5225_assgn52252 <= z5225_assgn52251;
        z5225_assgn52253 <= z5225_assgn52252;
        z1913_assgn1913 <= z5225_assgn52253;
        z5229_assgn52290 <= z5229_assgn5229;
        z5229_assgn52291 <= z5229_assgn52290;
        z5229_assgn52292 <= z5229_assgn52291;
        z5229_assgn52293 <= z5229_assgn52292;
        z1915_assgn1915 <= z5229_assgn52293;
        z5233_assgn52330 <= z5233_assgn5233;
        z5233_assgn52331 <= z5233_assgn52330;
        z5233_assgn52332 <= z5233_assgn52331;
        z5233_assgn52333 <= z5233_assgn52332;
        z1917_assgn1917 <= z5233_assgn52333;
        z5237_assgn52370 <= z5237_assgn5237;
        z5237_assgn52371 <= z5237_assgn52370;
        z5237_assgn52372 <= z5237_assgn52371;
        z5237_assgn52373 <= z5237_assgn52372;
        z1919_assgn1919 <= z5237_assgn52373;
        z5241_assgn52410 <= z5241_assgn5241;
        z5241_assgn52411 <= z5241_assgn52410;
        z5241_assgn52412 <= z5241_assgn52411;
        z5241_assgn52413 <= z5241_assgn52412;
        z1921_assgn1921 <= z5241_assgn52413;
        z5245_assgn52450 <= z5245_assgn5245;
        z5245_assgn52451 <= z5245_assgn52450;
        z5245_assgn52452 <= z5245_assgn52451;
        z5245_assgn52453 <= z5245_assgn52452;
        z1923_assgn1923 <= z5245_assgn52453;
        i1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg <= i1_hpc11_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc11_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc11_G4_mul1_G16_mul1_G256_inv0;
        i2_hpc11_G4_mul1_G16_mul1_G256_inv0_reg <= i2_hpc11_G4_mul1_G16_mul1_G256_inv0;
        p4_hpc11_G4_mul1_G16_mul1_G256_inv0_reg <= p4_hpc11_G4_mul1_G16_mul1_G256_inv0;
        z5265_assgn52650 <= z5265_assgn5265;
        z5265_assgn52651 <= z5265_assgn52650;
        z5265_assgn52652 <= z5265_assgn52651;
        z5265_assgn52653 <= z5265_assgn52652;
        z1941_assgn1941 <= z5265_assgn52653;
        z5269_assgn52690 <= z5269_assgn5269;
        z5269_assgn52691 <= z5269_assgn52690;
        z5269_assgn52692 <= z5269_assgn52691;
        z5269_assgn52693 <= z5269_assgn52692;
        z1943_assgn1943 <= z5269_assgn52693;
        z5273_assgn52730 <= z5273_assgn5273;
        z5273_assgn52731 <= z5273_assgn52730;
        z5273_assgn52732 <= z5273_assgn52731;
        z5273_assgn52733 <= z5273_assgn52732;
        z1945_assgn1945 <= z5273_assgn52733;
        z5277_assgn52770 <= z5277_assgn5277;
        z5277_assgn52771 <= z5277_assgn52770;
        z5277_assgn52772 <= z5277_assgn52771;
        z5277_assgn52773 <= z5277_assgn52772;
        z1947_assgn1947 <= z5277_assgn52773;
        z5281_assgn52810 <= z5281_assgn5281;
        z5281_assgn52811 <= z5281_assgn52810;
        z5281_assgn52812 <= z5281_assgn52811;
        z5281_assgn52813 <= z5281_assgn52812;
        z1949_assgn1949 <= z5281_assgn52813;
        z5285_assgn52850 <= z5285_assgn5285;
        z5285_assgn52851 <= z5285_assgn52850;
        z5285_assgn52852 <= z5285_assgn52851;
        z5285_assgn52853 <= z5285_assgn52852;
        z1951_assgn1951 <= z5285_assgn52853;
        i1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg <= i1_hpc12_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc12_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc12_G4_mul1_G16_mul1_G256_inv0;
        i2_hpc12_G4_mul1_G16_mul1_G256_inv0_reg <= i2_hpc12_G4_mul1_G16_mul1_G256_inv0;
        p4_hpc12_G4_mul1_G16_mul1_G256_inv0_reg <= p4_hpc12_G4_mul1_G16_mul1_G256_inv0;
        z5297_assgn52970 <= z5297_assgn5297;
        z5297_assgn52971 <= z5297_assgn52970;
        z5297_assgn52972 <= z5297_assgn52971;
        z5297_assgn52973 <= z5297_assgn52972;
        z5297_assgn52974 <= z5297_assgn52973;
        z1961_assgn1961 <= z5297_assgn52974;
        z5301_assgn53010 <= z5301_assgn5301;
        z5301_assgn53011 <= z5301_assgn53010;
        z5301_assgn53012 <= z5301_assgn53011;
        z5301_assgn53013 <= z5301_assgn53012;
        z5301_assgn53014 <= z5301_assgn53013;
        z1963_assgn1963 <= z5301_assgn53014;
        z5325_assgn53250 <= z5325_assgn5325;
        z5325_assgn53251 <= z5325_assgn53250;
        z5325_assgn53252 <= z5325_assgn53251;
        z5325_assgn53253 <= z5325_assgn53252;
        z1985_assgn1985 <= z5325_assgn53253;
        z5329_assgn53290 <= z5329_assgn5329;
        z5329_assgn53291 <= z5329_assgn53290;
        z5329_assgn53292 <= z5329_assgn53291;
        z5329_assgn53293 <= z5329_assgn53292;
        z1987_assgn1987 <= z5329_assgn53293;
        z5333_assgn53330 <= z5333_assgn5333;
        z5333_assgn53331 <= z5333_assgn53330;
        z5333_assgn53332 <= z5333_assgn53331;
        z5333_assgn53333 <= z5333_assgn53332;
        z1989_assgn1989 <= z5333_assgn53333;
        z5337_assgn53370 <= z5337_assgn5337;
        z5337_assgn53371 <= z5337_assgn53370;
        z5337_assgn53372 <= z5337_assgn53371;
        z5337_assgn53373 <= z5337_assgn53372;
        z1991_assgn1991 <= z5337_assgn53373;
        z5341_assgn53410 <= z5341_assgn5341;
        z5341_assgn53411 <= z5341_assgn53410;
        z5341_assgn53412 <= z5341_assgn53411;
        z5341_assgn53413 <= z5341_assgn53412;
        z1993_assgn1993 <= z5341_assgn53413;
        z5345_assgn53450 <= z5345_assgn5345;
        z5345_assgn53451 <= z5345_assgn53450;
        z5345_assgn53452 <= z5345_assgn53451;
        z5345_assgn53453 <= z5345_assgn53452;
        z1995_assgn1995 <= z5345_assgn53453;
        z5377_assgn53770 <= z5377_assgn5377;
        z5377_assgn53771 <= z5377_assgn53770;
        z5377_assgn53772 <= z5377_assgn53771;
        z5377_assgn53773 <= z5377_assgn53772;
        z2025_assgn2025 <= z5377_assgn53773;
        z5381_assgn53810 <= z5381_assgn5381;
        z5381_assgn53811 <= z5381_assgn53810;
        z5381_assgn53812 <= z5381_assgn53811;
        z5381_assgn53813 <= z5381_assgn53812;
        z2027_assgn2027 <= z5381_assgn53813;
        z5385_assgn53850 <= z5385_assgn5385;
        z5385_assgn53851 <= z5385_assgn53850;
        z5385_assgn53852 <= z5385_assgn53851;
        z5385_assgn53853 <= z5385_assgn53852;
        z2029_assgn2029 <= z5385_assgn53853;
        z5389_assgn53890 <= z5389_assgn5389;
        z5389_assgn53891 <= z5389_assgn53890;
        z5389_assgn53892 <= z5389_assgn53891;
        z5389_assgn53893 <= z5389_assgn53892;
        z2031_assgn2031 <= z5389_assgn53893;
        z5393_assgn53930 <= z5393_assgn5393;
        z5393_assgn53931 <= z5393_assgn53930;
        z5393_assgn53932 <= z5393_assgn53931;
        z5393_assgn53933 <= z5393_assgn53932;
        z2033_assgn2033 <= z5393_assgn53933;
        z5397_assgn53970 <= z5397_assgn5397;
        z5397_assgn53971 <= z5397_assgn53970;
        z5397_assgn53972 <= z5397_assgn53971;
        z5397_assgn53973 <= z5397_assgn53972;
        z2035_assgn2035 <= z5397_assgn53973;
        i1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg <= i1_hpc10_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc10_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc10_G4_mul2_G16_mul1_G256_inv0;
        i2_hpc10_G4_mul2_G16_mul1_G256_inv0_reg <= i2_hpc10_G4_mul2_G16_mul1_G256_inv0;
        p4_hpc10_G4_mul2_G16_mul1_G256_inv0_reg <= p4_hpc10_G4_mul2_G16_mul1_G256_inv0;
        z5413_assgn54130 <= z5413_assgn5413;
        z5413_assgn54131 <= z5413_assgn54130;
        z5413_assgn54132 <= z5413_assgn54131;
        z5413_assgn54133 <= z5413_assgn54132;
        z2049_assgn2049 <= z5413_assgn54133;
        z5417_assgn54170 <= z5417_assgn5417;
        z5417_assgn54171 <= z5417_assgn54170;
        z5417_assgn54172 <= z5417_assgn54171;
        z5417_assgn54173 <= z5417_assgn54172;
        z2051_assgn2051 <= z5417_assgn54173;
        z5421_assgn54210 <= z5421_assgn5421;
        z5421_assgn54211 <= z5421_assgn54210;
        z5421_assgn54212 <= z5421_assgn54211;
        z5421_assgn54213 <= z5421_assgn54212;
        z2053_assgn2053 <= z5421_assgn54213;
        z5425_assgn54250 <= z5425_assgn5425;
        z5425_assgn54251 <= z5425_assgn54250;
        z5425_assgn54252 <= z5425_assgn54251;
        z5425_assgn54253 <= z5425_assgn54252;
        z2055_assgn2055 <= z5425_assgn54253;
        z5429_assgn54290 <= z5429_assgn5429;
        z5429_assgn54291 <= z5429_assgn54290;
        z5429_assgn54292 <= z5429_assgn54291;
        z5429_assgn54293 <= z5429_assgn54292;
        z2057_assgn2057 <= z5429_assgn54293;
        z5433_assgn54330 <= z5433_assgn5433;
        z5433_assgn54331 <= z5433_assgn54330;
        z5433_assgn54332 <= z5433_assgn54331;
        z5433_assgn54333 <= z5433_assgn54332;
        z2059_assgn2059 <= z5433_assgn54333;
        i1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg <= i1_hpc11_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc11_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc11_G4_mul2_G16_mul1_G256_inv0;
        i2_hpc11_G4_mul2_G16_mul1_G256_inv0_reg <= i2_hpc11_G4_mul2_G16_mul1_G256_inv0;
        p4_hpc11_G4_mul2_G16_mul1_G256_inv0_reg <= p4_hpc11_G4_mul2_G16_mul1_G256_inv0;
        z5453_assgn54530 <= z5453_assgn5453;
        z5453_assgn54531 <= z5453_assgn54530;
        z5453_assgn54532 <= z5453_assgn54531;
        z5453_assgn54533 <= z5453_assgn54532;
        z2077_assgn2077 <= z5453_assgn54533;
        z5457_assgn54570 <= z5457_assgn5457;
        z5457_assgn54571 <= z5457_assgn54570;
        z5457_assgn54572 <= z5457_assgn54571;
        z5457_assgn54573 <= z5457_assgn54572;
        z2079_assgn2079 <= z5457_assgn54573;
        z5461_assgn54610 <= z5461_assgn5461;
        z5461_assgn54611 <= z5461_assgn54610;
        z5461_assgn54612 <= z5461_assgn54611;
        z5461_assgn54613 <= z5461_assgn54612;
        z2081_assgn2081 <= z5461_assgn54613;
        z5465_assgn54650 <= z5465_assgn5465;
        z5465_assgn54651 <= z5465_assgn54650;
        z5465_assgn54652 <= z5465_assgn54651;
        z5465_assgn54653 <= z5465_assgn54652;
        z2083_assgn2083 <= z5465_assgn54653;
        z5469_assgn54690 <= z5469_assgn5469;
        z5469_assgn54691 <= z5469_assgn54690;
        z5469_assgn54692 <= z5469_assgn54691;
        z5469_assgn54693 <= z5469_assgn54692;
        z2085_assgn2085 <= z5469_assgn54693;
        z5473_assgn54730 <= z5473_assgn5473;
        z5473_assgn54731 <= z5473_assgn54730;
        z5473_assgn54732 <= z5473_assgn54731;
        z5473_assgn54733 <= z5473_assgn54732;
        z2087_assgn2087 <= z5473_assgn54733;
        i1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg <= i1_hpc12_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc12_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc12_G4_mul2_G16_mul1_G256_inv0;
        i2_hpc12_G4_mul2_G16_mul1_G256_inv0_reg <= i2_hpc12_G4_mul2_G16_mul1_G256_inv0;
        p4_hpc12_G4_mul2_G16_mul1_G256_inv0_reg <= p4_hpc12_G4_mul2_G16_mul1_G256_inv0;
        z5485_assgn54850 <= z5485_assgn5485;
        z5485_assgn54851 <= z5485_assgn54850;
        z5485_assgn54852 <= z5485_assgn54851;
        z5485_assgn54853 <= z5485_assgn54852;
        z5485_assgn54854 <= z5485_assgn54853;
        z2097_assgn2097 <= z5485_assgn54854;
        z5489_assgn54890 <= z5489_assgn5489;
        z5489_assgn54891 <= z5489_assgn54890;
        z5489_assgn54892 <= z5489_assgn54891;
        z5489_assgn54893 <= z5489_assgn54892;
        z5489_assgn54894 <= z5489_assgn54893;
        z2099_assgn2099 <= z5489_assgn54894;
        z5501_assgn55010 <= z5501_assgn5501;
        z5501_assgn55011 <= z5501_assgn55010;
        z5501_assgn55012 <= z5501_assgn55011;
        z5501_assgn55013 <= z5501_assgn55012;
        z5501_assgn55014 <= z5501_assgn55013;
        z2109_assgn2109 <= z5501_assgn55014;
        z5505_assgn55050 <= z5505_assgn5505;
        z5505_assgn55051 <= z5505_assgn55050;
        z5505_assgn55052 <= z5505_assgn55051;
        z5505_assgn55053 <= z5505_assgn55052;
        z5505_assgn55054 <= z5505_assgn55053;
        z2111_assgn2111 <= z5505_assgn55054;
        z5549_assgn55490 <= z5549_assgn5549;
        z5549_assgn55491 <= z5549_assgn55490;
        z5549_assgn55492 <= z5549_assgn55491;
        z5549_assgn55493 <= z5549_assgn55492;
        z2153_assgn2153 <= z5549_assgn55493;
        z5553_assgn55530 <= z5553_assgn5553;
        z5553_assgn55531 <= z5553_assgn55530;
        z5553_assgn55532 <= z5553_assgn55531;
        z5553_assgn55533 <= z5553_assgn55532;
        z2155_assgn2155 <= z5553_assgn55533;
        z5557_assgn55570 <= z5557_assgn5557;
        z5557_assgn55571 <= z5557_assgn55570;
        z5557_assgn55572 <= z5557_assgn55571;
        z5557_assgn55573 <= z5557_assgn55572;
        z2157_assgn2157 <= z5557_assgn55573;
        z5561_assgn55610 <= z5561_assgn5561;
        z5561_assgn55611 <= z5561_assgn55610;
        z5561_assgn55612 <= z5561_assgn55611;
        z5561_assgn55613 <= z5561_assgn55612;
        z2159_assgn2159 <= z5561_assgn55613;
        z5565_assgn55650 <= z5565_assgn5565;
        z5565_assgn55651 <= z5565_assgn55650;
        z5565_assgn55652 <= z5565_assgn55651;
        z5565_assgn55653 <= z5565_assgn55652;
        z2161_assgn2161 <= z5565_assgn55653;
        z5569_assgn55690 <= z5569_assgn5569;
        z5569_assgn55691 <= z5569_assgn55690;
        z5569_assgn55692 <= z5569_assgn55691;
        z5569_assgn55693 <= z5569_assgn55692;
        z2163_assgn2163 <= z5569_assgn55693;
        z5605_assgn56050 <= z5605_assgn5605;
        z5605_assgn56051 <= z5605_assgn56050;
        z5605_assgn56052 <= z5605_assgn56051;
        z5605_assgn56053 <= z5605_assgn56052;
        z2197_assgn2197 <= z5605_assgn56053;
        z5609_assgn56090 <= z5609_assgn5609;
        z5609_assgn56091 <= z5609_assgn56090;
        z5609_assgn56092 <= z5609_assgn56091;
        z5609_assgn56093 <= z5609_assgn56092;
        z2199_assgn2199 <= z5609_assgn56093;
        z5613_assgn56130 <= z5613_assgn5613;
        z5613_assgn56131 <= z5613_assgn56130;
        z5613_assgn56132 <= z5613_assgn56131;
        z5613_assgn56133 <= z5613_assgn56132;
        z2201_assgn2201 <= z5613_assgn56133;
        z5617_assgn56170 <= z5617_assgn5617;
        z5617_assgn56171 <= z5617_assgn56170;
        z5617_assgn56172 <= z5617_assgn56171;
        z5617_assgn56173 <= z5617_assgn56172;
        z2203_assgn2203 <= z5617_assgn56173;
        z5621_assgn56210 <= z5621_assgn5621;
        z5621_assgn56211 <= z5621_assgn56210;
        z5621_assgn56212 <= z5621_assgn56211;
        z5621_assgn56213 <= z5621_assgn56212;
        z2205_assgn2205 <= z5621_assgn56213;
        z5625_assgn56250 <= z5625_assgn5625;
        z5625_assgn56251 <= z5625_assgn56250;
        z5625_assgn56252 <= z5625_assgn56251;
        z5625_assgn56253 <= z5625_assgn56252;
        z2207_assgn2207 <= z5625_assgn56253;
        z5657_assgn56570 <= z5657_assgn5657;
        z5657_assgn56571 <= z5657_assgn56570;
        z5657_assgn56572 <= z5657_assgn56571;
        z5657_assgn56573 <= z5657_assgn56572;
        z2237_assgn2237 <= z5657_assgn56573;
        z5661_assgn56610 <= z5661_assgn5661;
        z5661_assgn56611 <= z5661_assgn56610;
        z5661_assgn56612 <= z5661_assgn56611;
        z5661_assgn56613 <= z5661_assgn56612;
        z2239_assgn2239 <= z5661_assgn56613;
        z5665_assgn56650 <= z5665_assgn5665;
        z5665_assgn56651 <= z5665_assgn56650;
        z5665_assgn56652 <= z5665_assgn56651;
        z5665_assgn56653 <= z5665_assgn56652;
        z2241_assgn2241 <= z5665_assgn56653;
        z5669_assgn56690 <= z5669_assgn5669;
        z5669_assgn56691 <= z5669_assgn56690;
        z5669_assgn56692 <= z5669_assgn56691;
        z5669_assgn56693 <= z5669_assgn56692;
        z2243_assgn2243 <= z5669_assgn56693;
        z5673_assgn56730 <= z5673_assgn5673;
        z5673_assgn56731 <= z5673_assgn56730;
        z5673_assgn56732 <= z5673_assgn56731;
        z5673_assgn56733 <= z5673_assgn56732;
        z2245_assgn2245 <= z5673_assgn56733;
        z5677_assgn56770 <= z5677_assgn5677;
        z5677_assgn56771 <= z5677_assgn56770;
        z5677_assgn56772 <= z5677_assgn56771;
        z5677_assgn56773 <= z5677_assgn56772;
        z2247_assgn2247 <= z5677_assgn56773;
        i1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg <= i1_hpc10_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc10_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc10_G4_mul0_G16_mul2_G256_inv0;
        i2_hpc10_G4_mul0_G16_mul2_G256_inv0_reg <= i2_hpc10_G4_mul0_G16_mul2_G256_inv0;
        p4_hpc10_G4_mul0_G16_mul2_G256_inv0_reg <= p4_hpc10_G4_mul0_G16_mul2_G256_inv0;
        z5693_assgn56930 <= z5693_assgn5693;
        z5693_assgn56931 <= z5693_assgn56930;
        z5693_assgn56932 <= z5693_assgn56931;
        z5693_assgn56933 <= z5693_assgn56932;
        z2261_assgn2261 <= z5693_assgn56933;
        z5697_assgn56970 <= z5697_assgn5697;
        z5697_assgn56971 <= z5697_assgn56970;
        z5697_assgn56972 <= z5697_assgn56971;
        z5697_assgn56973 <= z5697_assgn56972;
        z2263_assgn2263 <= z5697_assgn56973;
        z5701_assgn57010 <= z5701_assgn5701;
        z5701_assgn57011 <= z5701_assgn57010;
        z5701_assgn57012 <= z5701_assgn57011;
        z5701_assgn57013 <= z5701_assgn57012;
        z2265_assgn2265 <= z5701_assgn57013;
        z5705_assgn57050 <= z5705_assgn5705;
        z5705_assgn57051 <= z5705_assgn57050;
        z5705_assgn57052 <= z5705_assgn57051;
        z5705_assgn57053 <= z5705_assgn57052;
        z2267_assgn2267 <= z5705_assgn57053;
        z5709_assgn57090 <= z5709_assgn5709;
        z5709_assgn57091 <= z5709_assgn57090;
        z5709_assgn57092 <= z5709_assgn57091;
        z5709_assgn57093 <= z5709_assgn57092;
        z2269_assgn2269 <= z5709_assgn57093;
        z5713_assgn57130 <= z5713_assgn5713;
        z5713_assgn57131 <= z5713_assgn57130;
        z5713_assgn57132 <= z5713_assgn57131;
        z5713_assgn57133 <= z5713_assgn57132;
        z2271_assgn2271 <= z5713_assgn57133;
        i1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg <= i1_hpc11_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc11_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc11_G4_mul0_G16_mul2_G256_inv0;
        i2_hpc11_G4_mul0_G16_mul2_G256_inv0_reg <= i2_hpc11_G4_mul0_G16_mul2_G256_inv0;
        p4_hpc11_G4_mul0_G16_mul2_G256_inv0_reg <= p4_hpc11_G4_mul0_G16_mul2_G256_inv0;
        z5733_assgn57330 <= z5733_assgn5733;
        z5733_assgn57331 <= z5733_assgn57330;
        z5733_assgn57332 <= z5733_assgn57331;
        z5733_assgn57333 <= z5733_assgn57332;
        z2289_assgn2289 <= z5733_assgn57333;
        z5737_assgn57370 <= z5737_assgn5737;
        z5737_assgn57371 <= z5737_assgn57370;
        z5737_assgn57372 <= z5737_assgn57371;
        z5737_assgn57373 <= z5737_assgn57372;
        z2291_assgn2291 <= z5737_assgn57373;
        z5741_assgn57410 <= z5741_assgn5741;
        z5741_assgn57411 <= z5741_assgn57410;
        z5741_assgn57412 <= z5741_assgn57411;
        z5741_assgn57413 <= z5741_assgn57412;
        z2293_assgn2293 <= z5741_assgn57413;
        z5745_assgn57450 <= z5745_assgn5745;
        z5745_assgn57451 <= z5745_assgn57450;
        z5745_assgn57452 <= z5745_assgn57451;
        z5745_assgn57453 <= z5745_assgn57452;
        z2295_assgn2295 <= z5745_assgn57453;
        z5749_assgn57490 <= z5749_assgn5749;
        z5749_assgn57491 <= z5749_assgn57490;
        z5749_assgn57492 <= z5749_assgn57491;
        z5749_assgn57493 <= z5749_assgn57492;
        z2297_assgn2297 <= z5749_assgn57493;
        z5753_assgn57530 <= z5753_assgn5753;
        z5753_assgn57531 <= z5753_assgn57530;
        z5753_assgn57532 <= z5753_assgn57531;
        z5753_assgn57533 <= z5753_assgn57532;
        z2299_assgn2299 <= z5753_assgn57533;
        i1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg <= i1_hpc12_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc12_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc12_G4_mul0_G16_mul2_G256_inv0;
        i2_hpc12_G4_mul0_G16_mul2_G256_inv0_reg <= i2_hpc12_G4_mul0_G16_mul2_G256_inv0;
        p4_hpc12_G4_mul0_G16_mul2_G256_inv0_reg <= p4_hpc12_G4_mul0_G16_mul2_G256_inv0;
        z5765_assgn57650 <= z5765_assgn5765;
        z5765_assgn57651 <= z5765_assgn57650;
        z5765_assgn57652 <= z5765_assgn57651;
        z5765_assgn57653 <= z5765_assgn57652;
        z5765_assgn57654 <= z5765_assgn57653;
        z2309_assgn2309 <= z5765_assgn57654;
        z5769_assgn57690 <= z5769_assgn5769;
        z5769_assgn57691 <= z5769_assgn57690;
        z5769_assgn57692 <= z5769_assgn57691;
        z5769_assgn57693 <= z5769_assgn57692;
        z5769_assgn57694 <= z5769_assgn57693;
        z2311_assgn2311 <= z5769_assgn57694;
        z5777_assgn57770 <= z5777_assgn5777;
        z5777_assgn57771 <= z5777_assgn57770;
        z5777_assgn57772 <= z5777_assgn57771;
        z5777_assgn57773 <= z5777_assgn57772;
        z5777_assgn57774 <= z5777_assgn57773;
        z2317_assgn2317 <= z5777_assgn57774;
        z5781_assgn57810 <= z5781_assgn5781;
        z5781_assgn57811 <= z5781_assgn57810;
        z5781_assgn57812 <= z5781_assgn57811;
        z5781_assgn57813 <= z5781_assgn57812;
        z5781_assgn57814 <= z5781_assgn57813;
        z2319_assgn2319 <= z5781_assgn57814;
        z5785_assgn57850 <= z5785_assgn5785;
        z5785_assgn57851 <= z5785_assgn57850;
        z5785_assgn57852 <= z5785_assgn57851;
        z5785_assgn57853 <= z5785_assgn57852;
        z5785_assgn57854 <= z5785_assgn57853;
        z2321_assgn2321 <= z5785_assgn57854;
        z5789_assgn57890 <= z5789_assgn5789;
        z5789_assgn57891 <= z5789_assgn57890;
        z5789_assgn57892 <= z5789_assgn57891;
        z5789_assgn57893 <= z5789_assgn57892;
        z5789_assgn57894 <= z5789_assgn57893;
        z2323_assgn2323 <= z5789_assgn57894;
        z5793_assgn57930 <= z5793_assgn5793;
        z5793_assgn57931 <= z5793_assgn57930;
        z5793_assgn57932 <= z5793_assgn57931;
        z5793_assgn57933 <= z5793_assgn57932;
        z5793_assgn57934 <= z5793_assgn57933;
        z2325_assgn2325 <= z5793_assgn57934;
        z5797_assgn57970 <= z5797_assgn5797;
        z5797_assgn57971 <= z5797_assgn57970;
        z5797_assgn57972 <= z5797_assgn57971;
        z5797_assgn57973 <= z5797_assgn57972;
        z5797_assgn57974 <= z5797_assgn57973;
        z2327_assgn2327 <= z5797_assgn57974;
        z5809_assgn58090 <= z5809_assgn5809;
        z5809_assgn58091 <= z5809_assgn58090;
        z5809_assgn58092 <= z5809_assgn58091;
        z5809_assgn58093 <= z5809_assgn58092;
        z5809_assgn58094 <= z5809_assgn58093;
        z2337_assgn2337 <= z5809_assgn58094;
        z5813_assgn58130 <= z5813_assgn5813;
        z5813_assgn58131 <= z5813_assgn58130;
        z5813_assgn58132 <= z5813_assgn58131;
        z5813_assgn58133 <= z5813_assgn58132;
        z5813_assgn58134 <= z5813_assgn58133;
        z2339_assgn2339 <= z5813_assgn58134;
        z5833_assgn58330 <= z5833_assgn5833;
        z5833_assgn58331 <= z5833_assgn58330;
        z5833_assgn58332 <= z5833_assgn58331;
        z5833_assgn58333 <= z5833_assgn58332;
        z2357_assgn2357 <= z5833_assgn58333;
        z5837_assgn58370 <= z5837_assgn5837;
        z5837_assgn58371 <= z5837_assgn58370;
        z5837_assgn58372 <= z5837_assgn58371;
        z5837_assgn58373 <= z5837_assgn58372;
        z2359_assgn2359 <= z5837_assgn58373;
        z5841_assgn58410 <= z5841_assgn5841;
        z5841_assgn58411 <= z5841_assgn58410;
        z5841_assgn58412 <= z5841_assgn58411;
        z5841_assgn58413 <= z5841_assgn58412;
        z2361_assgn2361 <= z5841_assgn58413;
        z5845_assgn58450 <= z5845_assgn5845;
        z5845_assgn58451 <= z5845_assgn58450;
        z5845_assgn58452 <= z5845_assgn58451;
        z5845_assgn58453 <= z5845_assgn58452;
        z2363_assgn2363 <= z5845_assgn58453;
        z5849_assgn58490 <= z5849_assgn5849;
        z5849_assgn58491 <= z5849_assgn58490;
        z5849_assgn58492 <= z5849_assgn58491;
        z5849_assgn58493 <= z5849_assgn58492;
        z2365_assgn2365 <= z5849_assgn58493;
        z5853_assgn58530 <= z5853_assgn5853;
        z5853_assgn58531 <= z5853_assgn58530;
        z5853_assgn58532 <= z5853_assgn58531;
        z5853_assgn58533 <= z5853_assgn58532;
        z2367_assgn2367 <= z5853_assgn58533;
        z5885_assgn58850 <= z5885_assgn5885;
        z5885_assgn58851 <= z5885_assgn58850;
        z5885_assgn58852 <= z5885_assgn58851;
        z5885_assgn58853 <= z5885_assgn58852;
        z2397_assgn2397 <= z5885_assgn58853;
        z5889_assgn58890 <= z5889_assgn5889;
        z5889_assgn58891 <= z5889_assgn58890;
        z5889_assgn58892 <= z5889_assgn58891;
        z5889_assgn58893 <= z5889_assgn58892;
        z2399_assgn2399 <= z5889_assgn58893;
        z5893_assgn58930 <= z5893_assgn5893;
        z5893_assgn58931 <= z5893_assgn58930;
        z5893_assgn58932 <= z5893_assgn58931;
        z5893_assgn58933 <= z5893_assgn58932;
        z2401_assgn2401 <= z5893_assgn58933;
        z5897_assgn58970 <= z5897_assgn5897;
        z5897_assgn58971 <= z5897_assgn58970;
        z5897_assgn58972 <= z5897_assgn58971;
        z5897_assgn58973 <= z5897_assgn58972;
        z2403_assgn2403 <= z5897_assgn58973;
        z5901_assgn59010 <= z5901_assgn5901;
        z5901_assgn59011 <= z5901_assgn59010;
        z5901_assgn59012 <= z5901_assgn59011;
        z5901_assgn59013 <= z5901_assgn59012;
        z2405_assgn2405 <= z5901_assgn59013;
        z5905_assgn59050 <= z5905_assgn5905;
        z5905_assgn59051 <= z5905_assgn59050;
        z5905_assgn59052 <= z5905_assgn59051;
        z5905_assgn59053 <= z5905_assgn59052;
        z2407_assgn2407 <= z5905_assgn59053;
        i1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg <= i1_hpc10_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc10_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc10_G4_mul1_G16_mul2_G256_inv0;
        i2_hpc10_G4_mul1_G16_mul2_G256_inv0_reg <= i2_hpc10_G4_mul1_G16_mul2_G256_inv0;
        p4_hpc10_G4_mul1_G16_mul2_G256_inv0_reg <= p4_hpc10_G4_mul1_G16_mul2_G256_inv0;
        z5921_assgn59210 <= z5921_assgn5921;
        z5921_assgn59211 <= z5921_assgn59210;
        z5921_assgn59212 <= z5921_assgn59211;
        z5921_assgn59213 <= z5921_assgn59212;
        z2421_assgn2421 <= z5921_assgn59213;
        z5925_assgn59250 <= z5925_assgn5925;
        z5925_assgn59251 <= z5925_assgn59250;
        z5925_assgn59252 <= z5925_assgn59251;
        z5925_assgn59253 <= z5925_assgn59252;
        z2423_assgn2423 <= z5925_assgn59253;
        z5929_assgn59290 <= z5929_assgn5929;
        z5929_assgn59291 <= z5929_assgn59290;
        z5929_assgn59292 <= z5929_assgn59291;
        z5929_assgn59293 <= z5929_assgn59292;
        z2425_assgn2425 <= z5929_assgn59293;
        z5933_assgn59330 <= z5933_assgn5933;
        z5933_assgn59331 <= z5933_assgn59330;
        z5933_assgn59332 <= z5933_assgn59331;
        z5933_assgn59333 <= z5933_assgn59332;
        z2427_assgn2427 <= z5933_assgn59333;
        z5937_assgn59370 <= z5937_assgn5937;
        z5937_assgn59371 <= z5937_assgn59370;
        z5937_assgn59372 <= z5937_assgn59371;
        z5937_assgn59373 <= z5937_assgn59372;
        z2429_assgn2429 <= z5937_assgn59373;
        z5941_assgn59410 <= z5941_assgn5941;
        z5941_assgn59411 <= z5941_assgn59410;
        z5941_assgn59412 <= z5941_assgn59411;
        z5941_assgn59413 <= z5941_assgn59412;
        z2431_assgn2431 <= z5941_assgn59413;
        i1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg <= i1_hpc11_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc11_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc11_G4_mul1_G16_mul2_G256_inv0;
        i2_hpc11_G4_mul1_G16_mul2_G256_inv0_reg <= i2_hpc11_G4_mul1_G16_mul2_G256_inv0;
        p4_hpc11_G4_mul1_G16_mul2_G256_inv0_reg <= p4_hpc11_G4_mul1_G16_mul2_G256_inv0;
        z5961_assgn59610 <= z5961_assgn5961;
        z5961_assgn59611 <= z5961_assgn59610;
        z5961_assgn59612 <= z5961_assgn59611;
        z5961_assgn59613 <= z5961_assgn59612;
        z2449_assgn2449 <= z5961_assgn59613;
        z5965_assgn59650 <= z5965_assgn5965;
        z5965_assgn59651 <= z5965_assgn59650;
        z5965_assgn59652 <= z5965_assgn59651;
        z5965_assgn59653 <= z5965_assgn59652;
        z2451_assgn2451 <= z5965_assgn59653;
        z5969_assgn59690 <= z5969_assgn5969;
        z5969_assgn59691 <= z5969_assgn59690;
        z5969_assgn59692 <= z5969_assgn59691;
        z5969_assgn59693 <= z5969_assgn59692;
        z2453_assgn2453 <= z5969_assgn59693;
        z5973_assgn59730 <= z5973_assgn5973;
        z5973_assgn59731 <= z5973_assgn59730;
        z5973_assgn59732 <= z5973_assgn59731;
        z5973_assgn59733 <= z5973_assgn59732;
        z2455_assgn2455 <= z5973_assgn59733;
        z5977_assgn59770 <= z5977_assgn5977;
        z5977_assgn59771 <= z5977_assgn59770;
        z5977_assgn59772 <= z5977_assgn59771;
        z5977_assgn59773 <= z5977_assgn59772;
        z2457_assgn2457 <= z5977_assgn59773;
        z5981_assgn59810 <= z5981_assgn5981;
        z5981_assgn59811 <= z5981_assgn59810;
        z5981_assgn59812 <= z5981_assgn59811;
        z5981_assgn59813 <= z5981_assgn59812;
        z2459_assgn2459 <= z5981_assgn59813;
        i1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg <= i1_hpc12_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc12_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc12_G4_mul1_G16_mul2_G256_inv0;
        i2_hpc12_G4_mul1_G16_mul2_G256_inv0_reg <= i2_hpc12_G4_mul1_G16_mul2_G256_inv0;
        p4_hpc12_G4_mul1_G16_mul2_G256_inv0_reg <= p4_hpc12_G4_mul1_G16_mul2_G256_inv0;
        z5993_assgn59930 <= z5993_assgn5993;
        z5993_assgn59931 <= z5993_assgn59930;
        z5993_assgn59932 <= z5993_assgn59931;
        z5993_assgn59933 <= z5993_assgn59932;
        z5993_assgn59934 <= z5993_assgn59933;
        z2469_assgn2469 <= z5993_assgn59934;
        z5997_assgn59970 <= z5997_assgn5997;
        z5997_assgn59971 <= z5997_assgn59970;
        z5997_assgn59972 <= z5997_assgn59971;
        z5997_assgn59973 <= z5997_assgn59972;
        z5997_assgn59974 <= z5997_assgn59973;
        z2471_assgn2471 <= z5997_assgn59974;
        z6021_assgn60210 <= z6021_assgn6021;
        z6021_assgn60211 <= z6021_assgn60210;
        z6021_assgn60212 <= z6021_assgn60211;
        z6021_assgn60213 <= z6021_assgn60212;
        z2493_assgn2493 <= z6021_assgn60213;
        z6025_assgn60250 <= z6025_assgn6025;
        z6025_assgn60251 <= z6025_assgn60250;
        z6025_assgn60252 <= z6025_assgn60251;
        z6025_assgn60253 <= z6025_assgn60252;
        z2495_assgn2495 <= z6025_assgn60253;
        z6029_assgn60290 <= z6029_assgn6029;
        z6029_assgn60291 <= z6029_assgn60290;
        z6029_assgn60292 <= z6029_assgn60291;
        z6029_assgn60293 <= z6029_assgn60292;
        z2497_assgn2497 <= z6029_assgn60293;
        z6033_assgn60330 <= z6033_assgn6033;
        z6033_assgn60331 <= z6033_assgn60330;
        z6033_assgn60332 <= z6033_assgn60331;
        z6033_assgn60333 <= z6033_assgn60332;
        z2499_assgn2499 <= z6033_assgn60333;
        z6037_assgn60370 <= z6037_assgn6037;
        z6037_assgn60371 <= z6037_assgn60370;
        z6037_assgn60372 <= z6037_assgn60371;
        z6037_assgn60373 <= z6037_assgn60372;
        z2501_assgn2501 <= z6037_assgn60373;
        z6041_assgn60410 <= z6041_assgn6041;
        z6041_assgn60411 <= z6041_assgn60410;
        z6041_assgn60412 <= z6041_assgn60411;
        z6041_assgn60413 <= z6041_assgn60412;
        z2503_assgn2503 <= z6041_assgn60413;
        z6073_assgn60730 <= z6073_assgn6073;
        z6073_assgn60731 <= z6073_assgn60730;
        z6073_assgn60732 <= z6073_assgn60731;
        z6073_assgn60733 <= z6073_assgn60732;
        z2533_assgn2533 <= z6073_assgn60733;
        z6077_assgn60770 <= z6077_assgn6077;
        z6077_assgn60771 <= z6077_assgn60770;
        z6077_assgn60772 <= z6077_assgn60771;
        z6077_assgn60773 <= z6077_assgn60772;
        z2535_assgn2535 <= z6077_assgn60773;
        z6081_assgn60810 <= z6081_assgn6081;
        z6081_assgn60811 <= z6081_assgn60810;
        z6081_assgn60812 <= z6081_assgn60811;
        z6081_assgn60813 <= z6081_assgn60812;
        z2537_assgn2537 <= z6081_assgn60813;
        z6085_assgn60850 <= z6085_assgn6085;
        z6085_assgn60851 <= z6085_assgn60850;
        z6085_assgn60852 <= z6085_assgn60851;
        z6085_assgn60853 <= z6085_assgn60852;
        z2539_assgn2539 <= z6085_assgn60853;
        z6089_assgn60890 <= z6089_assgn6089;
        z6089_assgn60891 <= z6089_assgn60890;
        z6089_assgn60892 <= z6089_assgn60891;
        z6089_assgn60893 <= z6089_assgn60892;
        z2541_assgn2541 <= z6089_assgn60893;
        z6093_assgn60930 <= z6093_assgn6093;
        z6093_assgn60931 <= z6093_assgn60930;
        z6093_assgn60932 <= z6093_assgn60931;
        z6093_assgn60933 <= z6093_assgn60932;
        z2543_assgn2543 <= z6093_assgn60933;
        i1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg <= i1_hpc10_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc10_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc10_G4_mul2_G16_mul2_G256_inv0;
        i2_hpc10_G4_mul2_G16_mul2_G256_inv0_reg <= i2_hpc10_G4_mul2_G16_mul2_G256_inv0;
        p4_hpc10_G4_mul2_G16_mul2_G256_inv0_reg <= p4_hpc10_G4_mul2_G16_mul2_G256_inv0;
        z6109_assgn61090 <= z6109_assgn6109;
        z6109_assgn61091 <= z6109_assgn61090;
        z6109_assgn61092 <= z6109_assgn61091;
        z6109_assgn61093 <= z6109_assgn61092;
        z2557_assgn2557 <= z6109_assgn61093;
        z6113_assgn61130 <= z6113_assgn6113;
        z6113_assgn61131 <= z6113_assgn61130;
        z6113_assgn61132 <= z6113_assgn61131;
        z6113_assgn61133 <= z6113_assgn61132;
        z2559_assgn2559 <= z6113_assgn61133;
        z6117_assgn61170 <= z6117_assgn6117;
        z6117_assgn61171 <= z6117_assgn61170;
        z6117_assgn61172 <= z6117_assgn61171;
        z6117_assgn61173 <= z6117_assgn61172;
        z2561_assgn2561 <= z6117_assgn61173;
        z6121_assgn61210 <= z6121_assgn6121;
        z6121_assgn61211 <= z6121_assgn61210;
        z6121_assgn61212 <= z6121_assgn61211;
        z6121_assgn61213 <= z6121_assgn61212;
        z2563_assgn2563 <= z6121_assgn61213;
        z6125_assgn61250 <= z6125_assgn6125;
        z6125_assgn61251 <= z6125_assgn61250;
        z6125_assgn61252 <= z6125_assgn61251;
        z6125_assgn61253 <= z6125_assgn61252;
        z2565_assgn2565 <= z6125_assgn61253;
        z6129_assgn61290 <= z6129_assgn6129;
        z6129_assgn61291 <= z6129_assgn61290;
        z6129_assgn61292 <= z6129_assgn61291;
        z6129_assgn61293 <= z6129_assgn61292;
        z2567_assgn2567 <= z6129_assgn61293;
        i1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg <= i1_hpc11_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc11_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc11_G4_mul2_G16_mul2_G256_inv0;
        i2_hpc11_G4_mul2_G16_mul2_G256_inv0_reg <= i2_hpc11_G4_mul2_G16_mul2_G256_inv0;
        p4_hpc11_G4_mul2_G16_mul2_G256_inv0_reg <= p4_hpc11_G4_mul2_G16_mul2_G256_inv0;
        z6149_assgn61490 <= z6149_assgn6149;
        z6149_assgn61491 <= z6149_assgn61490;
        z6149_assgn61492 <= z6149_assgn61491;
        z6149_assgn61493 <= z6149_assgn61492;
        z2585_assgn2585 <= z6149_assgn61493;
        z6153_assgn61530 <= z6153_assgn6153;
        z6153_assgn61531 <= z6153_assgn61530;
        z6153_assgn61532 <= z6153_assgn61531;
        z6153_assgn61533 <= z6153_assgn61532;
        z2587_assgn2587 <= z6153_assgn61533;
        z6157_assgn61570 <= z6157_assgn6157;
        z6157_assgn61571 <= z6157_assgn61570;
        z6157_assgn61572 <= z6157_assgn61571;
        z6157_assgn61573 <= z6157_assgn61572;
        z2589_assgn2589 <= z6157_assgn61573;
        z6161_assgn61610 <= z6161_assgn6161;
        z6161_assgn61611 <= z6161_assgn61610;
        z6161_assgn61612 <= z6161_assgn61611;
        z6161_assgn61613 <= z6161_assgn61612;
        z2591_assgn2591 <= z6161_assgn61613;
        z6165_assgn61650 <= z6165_assgn6165;
        z6165_assgn61651 <= z6165_assgn61650;
        z6165_assgn61652 <= z6165_assgn61651;
        z6165_assgn61653 <= z6165_assgn61652;
        z2593_assgn2593 <= z6165_assgn61653;
        z6169_assgn61690 <= z6169_assgn6169;
        z6169_assgn61691 <= z6169_assgn61690;
        z6169_assgn61692 <= z6169_assgn61691;
        z6169_assgn61693 <= z6169_assgn61692;
        z2595_assgn2595 <= z6169_assgn61693;
        i1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg <= i1_hpc12_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc12_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc12_G4_mul2_G16_mul2_G256_inv0;
        i2_hpc12_G4_mul2_G16_mul2_G256_inv0_reg <= i2_hpc12_G4_mul2_G16_mul2_G256_inv0;
        p4_hpc12_G4_mul2_G16_mul2_G256_inv0_reg <= p4_hpc12_G4_mul2_G16_mul2_G256_inv0;
        z6181_assgn61810 <= z6181_assgn6181;
        z6181_assgn61811 <= z6181_assgn61810;
        z6181_assgn61812 <= z6181_assgn61811;
        z6181_assgn61813 <= z6181_assgn61812;
        z6181_assgn61814 <= z6181_assgn61813;
        z2605_assgn2605 <= z6181_assgn61814;
        z6185_assgn61850 <= z6185_assgn6185;
        z6185_assgn61851 <= z6185_assgn61850;
        z6185_assgn61852 <= z6185_assgn61851;
        z6185_assgn61853 <= z6185_assgn61852;
        z6185_assgn61854 <= z6185_assgn61853;
        z2607_assgn2607 <= z6185_assgn61854;
        z6197_assgn61970 <= z6197_assgn6197;
        z6197_assgn61971 <= z6197_assgn61970;
        z6197_assgn61972 <= z6197_assgn61971;
        z6197_assgn61973 <= z6197_assgn61972;
        z6197_assgn61974 <= z6197_assgn61973;
        z2617_assgn2617 <= z6197_assgn61974;
        z6201_assgn62010 <= z6201_assgn6201;
        z6201_assgn62011 <= z6201_assgn62010;
        z6201_assgn62012 <= z6201_assgn62011;
        z6201_assgn62013 <= z6201_assgn62012;
        z6201_assgn62014 <= z6201_assgn62013;
        z2619_assgn2619 <= z6201_assgn62014;
        z6209_assgn62090 <= z6209_assgn6209;
        z6209_assgn62091 <= z6209_assgn62090;
        z6209_assgn62092 <= z6209_assgn62091;
        z6209_assgn62093 <= z6209_assgn62092;
        z6209_assgn62094 <= z6209_assgn62093;
        z2625_assgn2625 <= z6209_assgn62094;
        z6213_assgn62130 <= z6213_assgn6213;
        z6213_assgn62131 <= z6213_assgn62130;
        z6213_assgn62132 <= z6213_assgn62131;
        z6213_assgn62133 <= z6213_assgn62132;
        z6213_assgn62134 <= z6213_assgn62133;
        z2627_assgn2627 <= z6213_assgn62134;
        z6225_assgn62250 <= z6225_assgn6225;
        z6225_assgn62251 <= z6225_assgn62250;
        z6225_assgn62252 <= z6225_assgn62251;
        z6225_assgn62253 <= z6225_assgn62252;
        z6225_assgn62254 <= z6225_assgn62253;
        z2637_assgn2637 <= z6225_assgn62254;
        z6233_assgn62330 <= z6233_assgn6233;
        z6233_assgn62331 <= z6233_assgn62330;
        z6233_assgn62332 <= z6233_assgn62331;
        z6233_assgn62333 <= z6233_assgn62332;
        z6233_assgn62334 <= z6233_assgn62333;
        z2643_assgn2643 <= z6233_assgn62334;
        z6237_assgn62370 <= z6237_assgn6237;
        z6237_assgn62371 <= z6237_assgn62370;
        z6237_assgn62372 <= z6237_assgn62371;
        z6237_assgn62373 <= z6237_assgn62372;
        z6237_assgn62374 <= z6237_assgn62373;
        z2646_assgn2646 <= z6237_assgn62374;
        z6243_assgn62430 <= z6243_assgn6243;
        z6243_assgn62431 <= z6243_assgn62430;
        z6243_assgn62432 <= z6243_assgn62431;
        z6243_assgn62433 <= z6243_assgn62432;
        z6243_assgn62434 <= z6243_assgn62433;
        z2649_assgn2649 <= z6243_assgn62434;
        z6249_assgn62490 <= z6249_assgn6249;
        z6249_assgn62491 <= z6249_assgn62490;
        z6249_assgn62492 <= z6249_assgn62491;
        z6249_assgn62493 <= z6249_assgn62492;
        z6249_assgn62494 <= z6249_assgn62493;
        z2653_assgn2653 <= z6249_assgn62494;
        z6255_assgn62550 <= z6255_assgn6255;
        z6255_assgn62551 <= z6255_assgn62550;
        z6255_assgn62552 <= z6255_assgn62551;
        z6255_assgn62553 <= z6255_assgn62552;
        z6255_assgn62554 <= z6255_assgn62553;
        z2657_assgn2657 <= z6255_assgn62554;
        z6265_assgn62650 <= z6265_assgn6265;
        z6265_assgn62651 <= z6265_assgn62650;
        z6265_assgn62652 <= z6265_assgn62651;
        z6265_assgn62653 <= z6265_assgn62652;
        z6265_assgn62654 <= z6265_assgn62653;
        z2665_assgn2665 <= z6265_assgn62654;
        z6271_assgn62710 <= z6271_assgn6271;
        z6271_assgn62711 <= z6271_assgn62710;
        z6271_assgn62712 <= z6271_assgn62711;
        z6271_assgn62713 <= z6271_assgn62712;
        z6271_assgn62714 <= z6271_assgn62713;
        z2669_assgn2669 <= z6271_assgn62714;
        z6277_assgn62770 <= z6277_assgn6277;
        z6277_assgn62771 <= z6277_assgn62770;
        z6277_assgn62772 <= z6277_assgn62771;
        z6277_assgn62773 <= z6277_assgn62772;
        z6277_assgn62774 <= z6277_assgn62773;
        z2673_assgn2673 <= z6277_assgn62774;
        z6287_assgn62870 <= z6287_assgn6287;
        z6287_assgn62871 <= z6287_assgn62870;
        z6287_assgn62872 <= z6287_assgn62871;
        z6287_assgn62873 <= z6287_assgn62872;
        z6287_assgn62874 <= z6287_assgn62873;
        z2681_assgn2681 <= z6287_assgn62874;
        z6293_assgn62930 <= z6293_assgn6293;
        z6293_assgn62931 <= z6293_assgn62930;
        z6293_assgn62932 <= z6293_assgn62931;
        z6293_assgn62933 <= z6293_assgn62932;
        z6293_assgn62934 <= z6293_assgn62933;
        z2685_assgn2685 <= z6293_assgn62934;
        z6299_assgn62990 <= z6299_assgn6299;
        z6299_assgn62991 <= z6299_assgn62990;
        z6299_assgn62992 <= z6299_assgn62991;
        z6299_assgn62993 <= z6299_assgn62992;
        z6299_assgn62994 <= z6299_assgn62993;
        z2689_assgn2689 <= z6299_assgn62994;
        z6309_assgn63090 <= z6309_assgn6309;
        z6309_assgn63091 <= z6309_assgn63090;
        z6309_assgn63092 <= z6309_assgn63091;
        z6309_assgn63093 <= z6309_assgn63092;
        z6309_assgn63094 <= z6309_assgn63093;
        z2697_assgn2697 <= z6309_assgn63094;
        z6315_assgn63150 <= z6315_assgn6315;
        z6315_assgn63151 <= z6315_assgn63150;
        z6315_assgn63152 <= z6315_assgn63151;
        z6315_assgn63153 <= z6315_assgn63152;
        z6315_assgn63154 <= z6315_assgn63153;
        z2701_assgn2701 <= z6315_assgn63154;
        z6321_assgn63210 <= z6321_assgn6321;
        z6321_assgn63211 <= z6321_assgn63210;
        z6321_assgn63212 <= z6321_assgn63211;
        z6321_assgn63213 <= z6321_assgn63212;
        z6321_assgn63214 <= z6321_assgn63213;
        z2705_assgn2705 <= z6321_assgn63214;
        z6331_assgn63310 <= z6331_assgn6331;
        z6331_assgn63311 <= z6331_assgn63310;
        z6331_assgn63312 <= z6331_assgn63311;
        z6331_assgn63313 <= z6331_assgn63312;
        z6331_assgn63314 <= z6331_assgn63313;
        z2713_assgn2713 <= z6331_assgn63314;
        z6337_assgn63370 <= z6337_assgn6337;
        z6337_assgn63371 <= z6337_assgn63370;
        z6337_assgn63372 <= z6337_assgn63371;
        z6337_assgn63373 <= z6337_assgn63372;
        z6337_assgn63374 <= z6337_assgn63373;
        z2717_assgn2717 <= z6337_assgn63374;
        z6343_assgn63430 <= z6343_assgn6343;
        z6343_assgn63431 <= z6343_assgn63430;
        z6343_assgn63432 <= z6343_assgn63431;
        z6343_assgn63433 <= z6343_assgn63432;
        z6343_assgn63434 <= z6343_assgn63433;
        z2721_assgn2721 <= z6343_assgn63434;
        z6353_assgn63530 <= z6353_assgn6353;
        z6353_assgn63531 <= z6353_assgn63530;
        z6353_assgn63532 <= z6353_assgn63531;
        z6353_assgn63533 <= z6353_assgn63532;
        z6353_assgn63534 <= z6353_assgn63533;
        z2729_assgn2729 <= z6353_assgn63534;
        z6359_assgn63590 <= z6359_assgn6359;
        z6359_assgn63591 <= z6359_assgn63590;
        z6359_assgn63592 <= z6359_assgn63591;
        z6359_assgn63593 <= z6359_assgn63592;
        z6359_assgn63594 <= z6359_assgn63593;
        z2733_assgn2733 <= z6359_assgn63594;
        z6365_assgn63650 <= z6365_assgn6365;
        z6365_assgn63651 <= z6365_assgn63650;
        z6365_assgn63652 <= z6365_assgn63651;
        z6365_assgn63653 <= z6365_assgn63652;
        z6365_assgn63654 <= z6365_assgn63653;
        z2737_assgn2737 <= z6365_assgn63654;
        z6375_assgn63750 <= z6375_assgn6375;
        z6375_assgn63751 <= z6375_assgn63750;
        z6375_assgn63752 <= z6375_assgn63751;
        z6375_assgn63753 <= z6375_assgn63752;
        z6375_assgn63754 <= z6375_assgn63753;
        z2745_assgn2745 <= z6375_assgn63754;
        z6381_assgn63810 <= z6381_assgn6381;
        z6381_assgn63811 <= z6381_assgn63810;
        z6381_assgn63812 <= z6381_assgn63811;
        z6381_assgn63813 <= z6381_assgn63812;
        z6381_assgn63814 <= z6381_assgn63813;
        z2749_assgn2749 <= z6381_assgn63814;
        z6387_assgn63870 <= z6387_assgn6387;
        z6387_assgn63871 <= z6387_assgn63870;
        z6387_assgn63872 <= z6387_assgn63871;
        z6387_assgn63873 <= z6387_assgn63872;
        z6387_assgn63874 <= z6387_assgn63873;
        z2753_assgn2753 <= z6387_assgn63874;
        z6397_assgn63970 <= z6397_assgn6397;
        z6397_assgn63971 <= z6397_assgn63970;
        z6397_assgn63972 <= z6397_assgn63971;
        z6397_assgn63973 <= z6397_assgn63972;
        z6397_assgn63974 <= z6397_assgn63973;
        z2761_assgn2761 <= z6397_assgn63974;
        z6407_assgn64070 <= z6407_assgn6407;
        z6407_assgn64071 <= z6407_assgn64070;
        z6407_assgn64072 <= z6407_assgn64071;
        z6407_assgn64073 <= z6407_assgn64072;
        z6407_assgn64074 <= z6407_assgn64073;
        z2769_assgn2769 <= z6407_assgn64074;
        z6415_assgn64150 <= z6415_assgn6415;
        z6415_assgn64151 <= z6415_assgn64150;
        z6415_assgn64152 <= z6415_assgn64151;
        z6415_assgn64153 <= z6415_assgn64152;
        z6415_assgn64154 <= z6415_assgn64153;
        z2775_assgn2775 <= z6415_assgn64154;
        z6419_assgn64190 <= z6419_assgn6419;
        z6419_assgn64191 <= z6419_assgn64190;
        z6419_assgn64192 <= z6419_assgn64191;
        z6419_assgn64193 <= z6419_assgn64192;
        z6419_assgn64194 <= z6419_assgn64193;
        z2778_assgn2778 <= z6419_assgn64194;
        z6425_assgn64250 <= z6425_assgn6425;
        z6425_assgn64251 <= z6425_assgn64250;
        z6425_assgn64252 <= z6425_assgn64251;
        z6425_assgn64253 <= z6425_assgn64252;
        z6425_assgn64254 <= z6425_assgn64253;
        z2781_assgn2781 <= z6425_assgn64254;
        z6431_assgn64310 <= z6431_assgn6431;
        z6431_assgn64311 <= z6431_assgn64310;
        z6431_assgn64312 <= z6431_assgn64311;
        z6431_assgn64313 <= z6431_assgn64312;
        z6431_assgn64314 <= z6431_assgn64313;
        z2785_assgn2785 <= z6431_assgn64314;
        z6437_assgn64370 <= z6437_assgn6437;
        z6437_assgn64371 <= z6437_assgn64370;
        z6437_assgn64372 <= z6437_assgn64371;
        z6437_assgn64373 <= z6437_assgn64372;
        z6437_assgn64374 <= z6437_assgn64373;
        z2789_assgn2789 <= z6437_assgn64374;
        z6447_assgn64470 <= z6447_assgn6447;
        z6447_assgn64471 <= z6447_assgn64470;
        z6447_assgn64472 <= z6447_assgn64471;
        z6447_assgn64473 <= z6447_assgn64472;
        z6447_assgn64474 <= z6447_assgn64473;
        z2797_assgn2797 <= z6447_assgn64474;
        z6453_assgn64530 <= z6453_assgn6453;
        z6453_assgn64531 <= z6453_assgn64530;
        z6453_assgn64532 <= z6453_assgn64531;
        z6453_assgn64533 <= z6453_assgn64532;
        z6453_assgn64534 <= z6453_assgn64533;
        z2801_assgn2801 <= z6453_assgn64534;
        z6459_assgn64590 <= z6459_assgn6459;
        z6459_assgn64591 <= z6459_assgn64590;
        z6459_assgn64592 <= z6459_assgn64591;
        z6459_assgn64593 <= z6459_assgn64592;
        z6459_assgn64594 <= z6459_assgn64593;
        z2805_assgn2805 <= z6459_assgn64594;
        z6469_assgn64690 <= z6469_assgn6469;
        z6469_assgn64691 <= z6469_assgn64690;
        z6469_assgn64692 <= z6469_assgn64691;
        z6469_assgn64693 <= z6469_assgn64692;
        z6469_assgn64694 <= z6469_assgn64693;
        z2813_assgn2813 <= z6469_assgn64694;
        z6475_assgn64750 <= z6475_assgn6475;
        z6475_assgn64751 <= z6475_assgn64750;
        z6475_assgn64752 <= z6475_assgn64751;
        z6475_assgn64753 <= z6475_assgn64752;
        z6475_assgn64754 <= z6475_assgn64753;
        z2817_assgn2817 <= z6475_assgn64754;
        z6481_assgn64810 <= z6481_assgn6481;
        z6481_assgn64811 <= z6481_assgn64810;
        z6481_assgn64812 <= z6481_assgn64811;
        z6481_assgn64813 <= z6481_assgn64812;
        z6481_assgn64814 <= z6481_assgn64813;
        z2821_assgn2821 <= z6481_assgn64814;
        z6491_assgn64910 <= z6491_assgn6491;
        z6491_assgn64911 <= z6491_assgn64910;
        z6491_assgn64912 <= z6491_assgn64911;
        z6491_assgn64913 <= z6491_assgn64912;
        z6491_assgn64914 <= z6491_assgn64913;
        z2829_assgn2829 <= z6491_assgn64914;
        z6497_assgn64970 <= z6497_assgn6497;
        z6497_assgn64971 <= z6497_assgn64970;
        z6497_assgn64972 <= z6497_assgn64971;
        z6497_assgn64973 <= z6497_assgn64972;
        z6497_assgn64974 <= z6497_assgn64973;
        z2833_assgn2833 <= z6497_assgn64974;
        z6503_assgn65030 <= z6503_assgn6503;
        z6503_assgn65031 <= z6503_assgn65030;
        z6503_assgn65032 <= z6503_assgn65031;
        z6503_assgn65033 <= z6503_assgn65032;
        z6503_assgn65034 <= z6503_assgn65033;
        z2837_assgn2837 <= z6503_assgn65034;
        z6513_assgn65130 <= z6513_assgn6513;
        z6513_assgn65131 <= z6513_assgn65130;
        z6513_assgn65132 <= z6513_assgn65131;
        z6513_assgn65133 <= z6513_assgn65132;
        z6513_assgn65134 <= z6513_assgn65133;
        z2845_assgn2845 <= z6513_assgn65134;
        z6519_assgn65190 <= z6519_assgn6519;
        z6519_assgn65191 <= z6519_assgn65190;
        z6519_assgn65192 <= z6519_assgn65191;
        z6519_assgn65193 <= z6519_assgn65192;
        z6519_assgn65194 <= z6519_assgn65193;
        z2849_assgn2849 <= z6519_assgn65194;
        z6525_assgn65250 <= z6525_assgn6525;
        z6525_assgn65251 <= z6525_assgn65250;
        z6525_assgn65252 <= z6525_assgn65251;
        z6525_assgn65253 <= z6525_assgn65252;
        z6525_assgn65254 <= z6525_assgn65253;
        z2853_assgn2853 <= z6525_assgn65254;
        z6535_assgn65350 <= z6535_assgn6535;
        z6535_assgn65351 <= z6535_assgn65350;
        z6535_assgn65352 <= z6535_assgn65351;
        z6535_assgn65353 <= z6535_assgn65352;
        z6535_assgn65354 <= z6535_assgn65353;
        z2861_assgn2861 <= z6535_assgn65354;
        z6541_assgn65410 <= z6541_assgn6541;
        z6541_assgn65411 <= z6541_assgn65410;
        z6541_assgn65412 <= z6541_assgn65411;
        z6541_assgn65413 <= z6541_assgn65412;
        z6541_assgn65414 <= z6541_assgn65413;
        z2865_assgn2865 <= z6541_assgn65414;
        z6547_assgn65470 <= z6547_assgn6547;
        z6547_assgn65471 <= z6547_assgn65470;
        z6547_assgn65472 <= z6547_assgn65471;
        z6547_assgn65473 <= z6547_assgn65472;
        z6547_assgn65474 <= z6547_assgn65473;
        z2869_assgn2869 <= z6547_assgn65474;
        z6557_assgn65570 <= z6557_assgn6557;
        z6557_assgn65571 <= z6557_assgn65570;
        z6557_assgn65572 <= z6557_assgn65571;
        z6557_assgn65573 <= z6557_assgn65572;
        z6557_assgn65574 <= z6557_assgn65573;
        z2877_assgn2877 <= z6557_assgn65574;
        z6563_assgn65630 <= z6563_assgn6563;
        z6563_assgn65631 <= z6563_assgn65630;
        z6563_assgn65632 <= z6563_assgn65631;
        z6563_assgn65633 <= z6563_assgn65632;
        z6563_assgn65634 <= z6563_assgn65633;
        z2881_assgn2881 <= z6563_assgn65634;
        z6569_assgn65690 <= z6569_assgn6569;
        z6569_assgn65691 <= z6569_assgn65690;
        z6569_assgn65692 <= z6569_assgn65691;
        z6569_assgn65693 <= z6569_assgn65692;
        z6569_assgn65694 <= z6569_assgn65693;
        z2885_assgn2885 <= z6569_assgn65694;
        z6579_assgn65790 <= z6579_assgn6579;
        z6579_assgn65791 <= z6579_assgn65790;
        z6579_assgn65792 <= z6579_assgn65791;
        z6579_assgn65793 <= z6579_assgn65792;
        z6579_assgn65794 <= z6579_assgn65793;
        z2893_assgn2893 <= z6579_assgn65794;
        z6585_assgn65850 <= z6585_assgn6585;
        z6585_assgn65851 <= z6585_assgn65850;
        z6585_assgn65852 <= z6585_assgn65851;
        z6585_assgn65853 <= z6585_assgn65852;
        z6585_assgn65854 <= z6585_assgn65853;
        z2897_assgn2897 <= z6585_assgn65854;
        y0 <= (t6 ^ z2897_assgn2897);
        y1 <= t7;
    end

endmodule


        