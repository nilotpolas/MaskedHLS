module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    r6,
    r7,
    r8,
    r9,
    r10,
    r11,
    r12,
    r13,
    r14,
    r15,
    r16,
    r17,
    r18,
    r19,
    r20,
    r21,
    r22,
    r23,
    r24,
    r25,
    r26,
    r27,
    r28,
    r29,
    r30,
    r31,
    r32,
    r33,
    r34,
    r35,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1,
);
//INPUTS
    input [7:0] clk;
    input [7:0]  t0;
    input [7:0]  t1;
    input [7:0]  r0;
    input [7:0]  r1;
    input [7:0]  r2;
    input [7:0]  r3;
    input [7:0]  r4;
    input [7:0]  r5;
    input [7:0]  r6;
    input [7:0]  r7;
    input [7:0]  r8;
    input [7:0]  r9;
    input [7:0]  r10;
    input [7:0]  r11;
    input [7:0]  r12;
    input [7:0]  r13;
    input [7:0]  r14;
    input [7:0]  r15;
    input [7:0]  r16;
    input [7:0]  r17;
    input [7:0]  r18;
    input [7:0]  r19;
    input [7:0]  r20;
    input [7:0]  r21;
    input [7:0]  r22;
    input [7:0]  r23;
    input [7:0]  r24;
    input [7:0]  r25;
    input [7:0]  r26;
    input [7:0]  r27;
    input [7:0]  r28;
    input [7:0]  r29;
    input [7:0]  r30;
    input [7:0]  r31;
    input [7:0]  r32;
    input [7:0]  r33;
    input [7:0]  r34;
    input [7:0]  r35;
    input [7:0]  dec_0;
    input [7:0]  dec_1;
    input [7:0]  dec_255;
    input [7:0]  dec_169;
    input [7:0]  dec_129;
    input [7:0]  dec_9;
    input [7:0]  dec_72;
    input [7:0]  dec_242;
    input [7:0]  dec_243;
    input [7:0]  dec_152;
    input [7:0]  dec_240;
    input [7:0]  dec_4;
    input [7:0]  dec_15;
    input [7:0]  dec_12;
    input [7:0]  dec_2;
    input [7:0]  dec_3;
    input [7:0]  dec_16;
    input [7:0]  dec_36;
    input [7:0]  dec_220;
    input [7:0]  dec_11;
    input [7:0]  dec_158;
    input [7:0]  dec_45;
    input [7:0]  dec_88;
    input [7:0]  dec_99;
//OUTPUTS
    output reg [7:0]   y0;
    output reg [7:0]   y1;
//Intermediate values
    wire [7:0]  dec_99_inp;
    wire [7:0]  dec_88_inp;
    wire [7:0]  dec_45_inp;
    wire [7:0]  dec_158_inp;
    wire [7:0]  dec_11_inp;
    wire [7:0]  dec_220_inp;
    wire [7:0]  dec_36_inp;
    wire [7:0]  dec_16_inp;
    wire [7:0]  dec_3_inp;
    wire [7:0]  dec_2_inp;
    wire [7:0]  dec_12_inp;
    wire [7:0]  dec_15_inp;
    wire [7:0]  dec_4_inp;
    wire [7:0]  dec_240_inp;
    wire [7:0]  dec_152_inp;
    wire [7:0]  dec_243_inp;
    wire [7:0]  dec_242_inp;
    wire [7:0]  dec_72_inp;
    wire [7:0]  dec_9_inp;
    wire [7:0]  dec_129_inp;
    wire [7:0]  dec_169_inp;
    wire [7:0]  dec_255_inp;
    wire [7:0]  dec_1_inp;
    wire [7:0]  dec_0_inp;
    wire [7:0]  t0_inp;
    wire [7:0]  t1_inp;
    wire [7:0]  r0_inp;
    wire [7:0]  r1_inp;
    wire [7:0]  r2_inp;
    wire [7:0]  r3_inp;
    wire [7:0]  r4_inp;
    wire [7:0]  r5_inp;
    wire [7:0]  r6_inp;
    wire [7:0]  r7_inp;
    wire [7:0]  r8_inp;
    wire [7:0]  r9_inp;
    wire [7:0]  r10_inp;
    wire [7:0]  r11_inp;
    wire [7:0]  r12_inp;
    wire [7:0]  r13_inp;
    wire [7:0]  r14_inp;
    wire [7:0]  r15_inp;
    wire [7:0]  r16_inp;
    wire [7:0]  r17_inp;
    wire [7:0]  r18_inp;
    wire [7:0]  r19_inp;
    wire [7:0]  r20_inp;
    wire [7:0]  r21_inp;
    wire [7:0]  r22_inp;
    wire [7:0]  r23_inp;
    wire [7:0]  r24_inp;
    wire [7:0]  r25_inp;
    wire [7:0]  r26_inp;
    wire [7:0]  r27_inp;
    wire [7:0]  r28_inp;
    wire [7:0]  r29_inp;
    wire [7:0]  r30_inp;
    wire [7:0]  r31_inp;
    wire [7:0]  r32_inp;
    wire [7:0]  r33_inp;
    wire [7:0]  r34_inp;
    wire [7:0]  r35_inp;
    wire [7:0]  y_G256_newbasis0;
    wire [7:0]  tempy1_G256_newbasis0;
    wire [7:0]  cond1_G256_newbasis0;
    wire [7:0]  negCond1_G256_newbasis0;
    wire [7:0]  yxorb1_G256_newbasis0;
    wire [7:0]  ny1_G256_newbasis0;
    wire [7:0]  tempybooloNegCond1_G256_newbasis0;
    wire [7:0]  y1_G256_newbasis0;
    wire [7:0]  x1_G256_newbasis0;
    wire [7:0]  tempy2_G256_newbasis0;
    wire [7:0]  cond2_G256_newbasis0;
    wire [7:0]  negCond2_G256_newbasis0;
    wire [7:0]  yxorb2_G256_newbasis0;
    wire [7:0]  ny2_G256_newbasis0;
    wire [7:0]  tempybooloNegCond2_G256_newbasis0;
    wire [7:0]  y2_G256_newbasis0;
    wire [7:0]  x2_G256_newbasis0;
    wire [7:0]  tempy3_G256_newbasis0;
    wire [7:0]  cond3_G256_newbasis0;
    wire [7:0]  negCond3_G256_newbasis0;
    wire [7:0]  yxorb3_G256_newbasis0;
    wire [7:0]  ny3_G256_newbasis0;
    wire [7:0]  tempybooloNegCond3_G256_newbasis0;
    wire [7:0]  y3_G256_newbasis0;
    wire [7:0]  x3_G256_newbasis0;
    wire [7:0]  tempy4_G256_newbasis0;
    wire [7:0]  cond4_G256_newbasis0;
    wire [7:0]  negCond4_G256_newbasis0;
    wire [7:0]  yxorb4_G256_newbasis0;
    wire [7:0]  ny4_G256_newbasis0;
    wire [7:0]  tempybooloNegCond4_G256_newbasis0;
    wire [7:0]  y4_G256_newbasis0;
    wire [7:0]  x4_G256_newbasis0;
    wire [7:0]  tempy5_G256_newbasis0;
    wire [7:0]  cond5_G256_newbasis0;
    wire [7:0]  negCond5_G256_newbasis0;
    wire [7:0]  yxorb5_G256_newbasis0;
    wire [7:0]  ny5_G256_newbasis0;
    wire [7:0]  tempybooloNegCond5_G256_newbasis0;
    wire [7:0]  y5_G256_newbasis0;
    wire [7:0]  x5_G256_newbasis0;
    wire [7:0]  tempy6_G256_newbasis0;
    wire [7:0]  cond6_G256_newbasis0;
    wire [7:0]  negCond6_G256_newbasis0;
    wire [7:0]  yxorb6_G256_newbasis0;
    wire [7:0]  ny6_G256_newbasis0;
    wire [7:0]  tempybooloNegCond6_G256_newbasis0;
    wire [7:0]  y6_G256_newbasis0;
    wire [7:0]  x6_G256_newbasis0;
    wire [7:0]  tempy7_G256_newbasis0;
    wire [7:0]  cond7_G256_newbasis0;
    wire [7:0]  negCond7_G256_newbasis0;
    wire [7:0]  yxorb7_G256_newbasis0;
    wire [7:0]  ny7_G256_newbasis0;
    wire [7:0]  tempybooloNegCond7_G256_newbasis0;
    wire [7:0]  y7_G256_newbasis0;
    wire [7:0]  x7_G256_newbasis0;
    wire [7:0]  tempy8_G256_newbasis0;
    wire [7:0]  cond8_G256_newbasis0;
    wire [7:0]  negCond8_G256_newbasis0;
    wire [7:0]  yxorb8_G256_newbasis0;
    wire [7:0]  ny8_G256_newbasis0;
    wire [7:0]  tempybooloNegCond8_G256_newbasis0;
    wire [7:0]  y8_G256_newbasis0;
    wire [7:0]  z2721_assgn2721;
    reg [7:0]  z2721_assgn27210;
    reg [7:0]  z2721_assgn27211;
    reg [7:0]  z2721_assgn27212;
    reg [7:0]  x8_G256_newbasis0;
    wire [7:0]  t2;
    wire [7:0]  z_y_G256_newbasis0;
    wire [7:0]  z_tempy1_G256_newbasis0;
    wire [7:0]  z_cond1_G256_newbasis0;
    wire [7:0]  z_negCond1_G256_newbasis0;
    wire [7:0]  z_yxorb1_G256_newbasis0;
    wire [7:0]  z_ny1_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond1_G256_newbasis0;
    wire [7:0]  z_y1_G256_newbasis0;
    wire [7:0]  z_x1_G256_newbasis0;
    wire [7:0]  z_tempy2_G256_newbasis0;
    wire [7:0]  z_cond2_G256_newbasis0;
    wire [7:0]  z_negCond2_G256_newbasis0;
    wire [7:0]  z_yxorb2_G256_newbasis0;
    wire [7:0]  z_ny2_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond2_G256_newbasis0;
    wire [7:0]  z_y2_G256_newbasis0;
    wire [7:0]  z_x2_G256_newbasis0;
    wire [7:0]  z_tempy3_G256_newbasis0;
    wire [7:0]  z_cond3_G256_newbasis0;
    wire [7:0]  z_negCond3_G256_newbasis0;
    wire [7:0]  z_yxorb3_G256_newbasis0;
    wire [7:0]  z_ny3_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond3_G256_newbasis0;
    wire [7:0]  z_y3_G256_newbasis0;
    wire [7:0]  z_x3_G256_newbasis0;
    wire [7:0]  z_tempy4_G256_newbasis0;
    wire [7:0]  z_cond4_G256_newbasis0;
    wire [7:0]  z_negCond4_G256_newbasis0;
    wire [7:0]  z_yxorb4_G256_newbasis0;
    wire [7:0]  z_ny4_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond4_G256_newbasis0;
    wire [7:0]  z_y4_G256_newbasis0;
    wire [7:0]  z_x4_G256_newbasis0;
    wire [7:0]  z_tempy5_G256_newbasis0;
    wire [7:0]  z_cond5_G256_newbasis0;
    wire [7:0]  z_negCond5_G256_newbasis0;
    wire [7:0]  z_yxorb5_G256_newbasis0;
    wire [7:0]  z_ny5_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond5_G256_newbasis0;
    wire [7:0]  z_y5_G256_newbasis0;
    wire [7:0]  z_x5_G256_newbasis0;
    wire [7:0]  z_tempy6_G256_newbasis0;
    wire [7:0]  z_cond6_G256_newbasis0;
    wire [7:0]  z_negCond6_G256_newbasis0;
    wire [7:0]  z_yxorb6_G256_newbasis0;
    wire [7:0]  z_ny6_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond6_G256_newbasis0;
    wire [7:0]  z_y6_G256_newbasis0;
    wire [7:0]  z_x6_G256_newbasis0;
    wire [7:0]  z_tempy7_G256_newbasis0;
    wire [7:0]  z_cond7_G256_newbasis0;
    wire [7:0]  z_negCond7_G256_newbasis0;
    wire [7:0]  z_yxorb7_G256_newbasis0;
    wire [7:0]  z_ny7_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond7_G256_newbasis0;
    wire [7:0]  z_y7_G256_newbasis0;
    wire [7:0]  z_x7_G256_newbasis0;
    wire [7:0]  z_tempy8_G256_newbasis0;
    wire [7:0]  z_cond8_G256_newbasis0;
    wire [7:0]  z_negCond8_G256_newbasis0;
    wire [7:0]  z_yxorb8_G256_newbasis0;
    wire [7:0]  z_ny8_G256_newbasis0;
    wire [7:0]  z_tempybooloNegCond8_G256_newbasis0;
    wire [7:0]  z_y8_G256_newbasis0;
    wire [7:0]  z2853_assgn2853;
    reg [7:0]  z2853_assgn28530;
    reg [7:0]  z2853_assgn28531;
    reg [7:0]  z2853_assgn28532;
    reg [7:0]  z_x8_G256_newbasis0;
    wire [7:0]  t3;
    wire [7:0]  a0_0_G256_inv0;
    wire [7:0]  a1_0_G256_inv0;
    wire [7:0]  a0_G256_inv0;
    wire [7:0]  a1_G256_inv0;
    wire [7:0]  b0_G256_inv0;
    wire [7:0]  b1_G256_inv0;
    wire [7:0]  a0xorb0_G256_inv0;
    wire [7:0]  a1xorb1_G256_inv0;
    wire [7:0]  a0_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1_G16_sq_scl0_G256_inv0;
    wire [7:0]  p0_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  p1_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0]  p0_G16_sq_scl0_G256_inv0;
    wire [7:0]  p1_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0]  q0_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  q1_0_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0]  q0_G16_sq_scl0_G256_inv0;
    wire [7:0]  q1_G16_sq_scl0_G256_inv0;
    wire [7:0]  p0ls2_G16_sq_scl0_G256_inv0;
    wire [7:0]  p1ls2_G16_sq_scl0_G256_inv0;
    wire [7:0]  c0_G256_inv0;
    wire [7:0]  c1_G256_inv0;
    wire [7:0]  r00_G16_mul0_G256_inv0;
    wire [7:0]  r10_G16_mul0_G256_inv0;
    wire [7:0]  r20_G16_mul0_G256_inv0;
    wire [7:0]  r30_G16_mul0_G256_inv0;
    wire [7:0]  r40_G16_mul0_G256_inv0;
    wire [7:0]  r50_G16_mul0_G256_inv0;
    wire [7:0]  r60_G16_mul0_G256_inv0;
    wire [7:0]  r70_G16_mul0_G256_inv0;
    wire [7:0]  r80_G16_mul0_G256_inv0;
    wire [7:0]  a0_0_G16_mul0_G256_inv0;
    wire [7:0]  a1_0_G16_mul0_G256_inv0;
    wire [7:0]  a0_G16_mul0_G256_inv0;
    wire [7:0]  a1_G16_mul0_G256_inv0;
    wire [7:0]  b0_G16_mul0_G256_inv0;
    wire [7:0]  b1_G16_mul0_G256_inv0;
    wire [7:0]  c0_0_G16_mul0_G256_inv0;
    wire [7:0]  c1_0_G16_mul0_G256_inv0;
    wire [7:0]  c0_G16_mul0_G256_inv0;
    wire [7:0]  c1_G16_mul0_G256_inv0;
    wire [7:0]  d0_G16_mul0_G256_inv0;
    wire [7:0]  d1_G16_mul0_G256_inv0;
    wire [7:0]  axorb_0_G16_mul0_G256_inv0;
    wire [7:0]  cxord_0_G16_mul0_G256_inv0;
    wire [7:0]  axorb_1_G16_mul0_G256_inv0;
    wire [7:0]  cxord_1_G16_mul0_G256_inv0;
    wire [7:0]  r00_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  r10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  r20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  a0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  a1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  b0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  b1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  c0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  c1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  d0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  d1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  q0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  q1_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0]  dec_1_inp_reg;
    wire [7:0]  p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0]  e0_G16_mul0_G256_inv0;
    wire [7:0]  e1_G16_mul0_G256_inv0;
    reg [7:0]  dec_2_inp_reg;
    wire [7:0]  a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0]  e01_G16_mul0_G256_inv0;
    wire [7:0]  e11_G16_mul0_G256_inv0;
    wire [7:0]  r00_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  r10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  r20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  a0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  a1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  b0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  b1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  c0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  c1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  d0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  d1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  q0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  q1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0]  p0_0_G16_mul0_G256_inv0;
    wire [7:0]  p1_0_G16_mul0_G256_inv0;
    wire [7:0]  p0_G16_mul0_G256_inv0;
    wire [7:0]  p1_G16_mul0_G256_inv0;
    wire [7:0]  r00_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  r10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  r20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  a0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  a1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  b0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  b1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  c0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  c1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  d0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  d1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p2_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i1_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p3_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  i2_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  q0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  q1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0]  q0_0_G16_mul0_G256_inv0;
    wire [7:0]  q1_0_G16_mul0_G256_inv0;
    wire [7:0]  q0_G16_mul0_G256_inv0;
    wire [7:0]  q1_G16_mul0_G256_inv0;
    wire [7:0]  p0ls2_G16_mul0_G256_inv0;
    wire [7:0]  p1ls2_G16_mul0_G256_inv0;
    wire [7:0]  d0_G256_inv0;
    wire [7:0]  d1_G256_inv0;
    reg [7:0]  c0_G256_inv0_reg;
    wire [7:0]  c0xord0_G256_inv0;
    reg [7:0]  c1_G256_inv0_reg;
    wire [7:0]  c1xord1_G256_inv0;
    wire [7:0]  r00_G16_inv0_G256_inv0;
    wire [7:0]  r10_G16_inv0_G256_inv0;
    wire [7:0]  r20_G16_inv0_G256_inv0;
    wire [7:0]  r30_G16_inv0_G256_inv0;
    wire [7:0]  r40_G16_inv0_G256_inv0;
    wire [7:0]  r50_G16_inv0_G256_inv0;
    wire [7:0]  r60_G16_inv0_G256_inv0;
    wire [7:0]  r70_G16_inv0_G256_inv0;
    wire [7:0]  r80_G16_inv0_G256_inv0;
    reg [7:0]  dec_12_inp_reg;
    wire [7:0]  a0_0_G16_inv0_G256_inv0;
    wire [7:0]  a1_0_G16_inv0_G256_inv0;
    wire [7:0]  a0_G16_inv0_G256_inv0;
    wire [7:0]  a1_G16_inv0_G256_inv0;
    reg [7:0]  dec_3_inp_reg;
    wire [7:0]  b0_G16_inv0_G256_inv0;
    wire [7:0]  b1_G16_inv0_G256_inv0;
    wire [7:0]  a0xorb0_G16_inv0_G256_inv0;
    wire [7:0]  a1xorb1_G16_inv0_G256_inv0;
    wire [7:0]  a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  a0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  a1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  b0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  b1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0]  c0_0_G16_inv0_G256_inv0;
    wire [7:0]  c1_0_G16_inv0_G256_inv0;
    wire [7:0]  a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0]  c0_G16_inv0_G256_inv0;
    wire [7:0]  c1_G16_inv0_G256_inv0;
    wire [7:0]  r00_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  r10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  r20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  a0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  a1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  b0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  b1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  c0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  c1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  d0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  d1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p2_domand0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  z0_domand0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  i1_domand0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p3_domand0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  i2_domand0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p2_domand1_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  z0_domand1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  i1_domand1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p3_domand1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  i2_domand1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p2_domand2_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  z0_domand2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  i1_domand2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p3_domand2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  i2_domand2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  q0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  q1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  z3569_assgn3569;
    reg [7:0]  z3569_assgn35690;
    reg [7:0]  z1101_assgn1101;
    wire [7:0]  p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  z3573_assgn3573;
    reg [7:0]  z3573_assgn35730;
    reg [7:0]  z1103_assgn1103;
    wire [7:0]  p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0]  d0_G16_inv0_G256_inv0;
    wire [7:0]  d1_G16_inv0_G256_inv0;
    reg [7:0]  c0_G16_inv0_G256_inv0_reg;
    wire [7:0]  c0xord0_G16_inv0_G256_inv0;
    reg [7:0]  c1_G16_inv0_G256_inv0_reg;
    wire [7:0]  c1xord1_G16_inv0_G256_inv0;
    wire [7:0]  z3585_assgn3585;
    reg [7:0]  z3585_assgn35850;
    reg [7:0]  z1113_assgn1113;
    wire [7:0]  a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3589_assgn3589;
    reg [7:0]  z3589_assgn35890;
    reg [7:0]  z1115_assgn1115;
    wire [7:0]  a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3593_assgn3593;
    reg [7:0]  z3593_assgn35930;
    reg [7:0]  z1117_assgn1117;
    wire [7:0]  a0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3597_assgn3597;
    reg [7:0]  z3597_assgn35970;
    reg [7:0]  z1119_assgn1119;
    wire [7:0]  a1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3601_assgn3601;
    reg [7:0]  z3601_assgn36010;
    reg [7:0]  z1121_assgn1121;
    wire [7:0]  b0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3605_assgn3605;
    reg [7:0]  z3605_assgn36050;
    reg [7:0]  z1123_assgn1123;
    wire [7:0]  b1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3609_assgn3609;
    reg [7:0]  z3609_assgn36090;
    reg [7:0]  z1125_assgn1125;
    wire [7:0]  b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  z3613_assgn3613;
    reg [7:0]  z3613_assgn36130;
    reg [7:0]  z1127_assgn1127;
    wire [7:0]  b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0]  e0_G16_inv0_G256_inv0;
    wire [7:0]  e1_G16_inv0_G256_inv0;
    wire [7:0]  r00_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  r10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  r20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3627_assgn3627;
    reg [7:0]  z3627_assgn36270;
    reg [7:0]  z1139_assgn1139;
    wire [7:0]  a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3631_assgn3631;
    reg [7:0]  z3631_assgn36310;
    reg [7:0]  z1141_assgn1141;
    wire [7:0]  a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3635_assgn3635;
    reg [7:0]  z3635_assgn36350;
    reg [7:0]  z1143_assgn1143;
    wire [7:0]  a0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3639_assgn3639;
    reg [7:0]  z3639_assgn36390;
    reg [7:0]  z1145_assgn1145;
    wire [7:0]  a1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3643_assgn3643;
    reg [7:0]  z3643_assgn36430;
    reg [7:0]  z1147_assgn1147;
    wire [7:0]  b0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3647_assgn3647;
    reg [7:0]  z3647_assgn36470;
    reg [7:0]  z1149_assgn1149;
    wire [7:0]  b1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  c0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  c1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  d0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  d1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  cxord_1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3675_assgn3675;
    reg [7:0]  z3675_assgn36750;
    reg [7:0]  z1175_assgn1175;
    wire [7:0]  i1_domand0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  cxord_0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3681_assgn3681;
    reg [7:0]  z3681_assgn36810;
    reg [7:0]  z1179_assgn1179;
    wire [7:0]  i2_domand0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  c1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3697_assgn3697;
    reg [7:0]  z3697_assgn36970;
    reg [7:0]  z1193_assgn1193;
    wire [7:0]  i1_domand1_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  c0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3703_assgn3703;
    reg [7:0]  z3703_assgn37030;
    reg [7:0]  z1197_assgn1197;
    wire [7:0]  i2_domand1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  d1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3723_assgn3723;
    reg [7:0]  z3723_assgn37230;
    reg [7:0]  z1215_assgn1215;
    wire [7:0]  i1_domand2_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  d0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3729_assgn3729;
    reg [7:0]  z3729_assgn37290;
    reg [7:0]  z1219_assgn1219;
    wire [7:0]  i2_domand2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  q0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  q1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3745_assgn3745;
    reg [7:0]  z3745_assgn37450;
    reg [7:0]  z3745_assgn37451;
    reg [7:0]  z1233_assgn1233;
    wire [7:0]  p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  z3749_assgn3749;
    reg [7:0]  z3749_assgn37490;
    reg [7:0]  z3749_assgn37491;
    reg [7:0]  z1235_assgn1235;
    wire [7:0]  p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0]  p0_G16_inv0_G256_inv0;
    wire [7:0]  p1_G16_inv0_G256_inv0;
    wire [7:0]  r00_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  r10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  r20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3763_assgn3763;
    reg [7:0]  z3763_assgn37630;
    reg [7:0]  z1247_assgn1247;
    wire [7:0]  a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3767_assgn3767;
    reg [7:0]  z3767_assgn37670;
    reg [7:0]  z1249_assgn1249;
    wire [7:0]  a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3771_assgn3771;
    reg [7:0]  z3771_assgn37710;
    reg [7:0]  z1251_assgn1251;
    wire [7:0]  a0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3775_assgn3775;
    reg [7:0]  z3775_assgn37750;
    reg [7:0]  z1253_assgn1253;
    wire [7:0]  a1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3779_assgn3779;
    reg [7:0]  z3779_assgn37790;
    reg [7:0]  z1255_assgn1255;
    wire [7:0]  b0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3783_assgn3783;
    reg [7:0]  z3783_assgn37830;
    reg [7:0]  z1257_assgn1257;
    wire [7:0]  b1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  c0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  c1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  d0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  d1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  axorb_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  cxord_1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3811_assgn3811;
    reg [7:0]  z3811_assgn38110;
    reg [7:0]  z1283_assgn1283;
    wire [7:0]  i1_domand0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  cxord_0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3817_assgn3817;
    reg [7:0]  z3817_assgn38170;
    reg [7:0]  z1287_assgn1287;
    wire [7:0]  i2_domand0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand0_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  e0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand0_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  e1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  c1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3833_assgn3833;
    reg [7:0]  z3833_assgn38330;
    reg [7:0]  z1301_assgn1301;
    wire [7:0]  i1_domand1_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  c0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3839_assgn3839;
    reg [7:0]  z3839_assgn38390;
    reg [7:0]  z1305_assgn1305;
    wire [7:0]  i2_domand1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand1_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand1_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand1_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  d1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p2_domand2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3859_assgn3859;
    reg [7:0]  z3859_assgn38590;
    reg [7:0]  z1323_assgn1323;
    wire [7:0]  i1_domand2_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  d0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  p3_domand2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3865_assgn3865;
    reg [7:0]  z3865_assgn38650;
    reg [7:0]  z1327_assgn1327;
    wire [7:0]  i2_domand2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p1_domand2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  p4_domand2_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i1_domand2_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p1_domand2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0]  i2_domand2_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0]  p4_domand2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  q0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  q1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3881_assgn3881;
    reg [7:0]  z3881_assgn38810;
    reg [7:0]  z3881_assgn38811;
    reg [7:0]  z1341_assgn1341;
    wire [7:0]  p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  z3885_assgn3885;
    reg [7:0]  z3885_assgn38850;
    reg [7:0]  z3885_assgn38851;
    reg [7:0]  z1343_assgn1343;
    wire [7:0]  p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0]  q0_G16_inv0_G256_inv0;
    wire [7:0]  q1_G16_inv0_G256_inv0;
    wire [7:0]  z3893_assgn3893;
    reg [7:0]  z3893_assgn38930;
    reg [7:0] z3893_assgn38931;
    reg [7:0] z1349_assgn1349;
    wire [7:0]  p0ls2_G16_inv0_G256_inv0;
    wire [7:0]  z3897_assgn3897;
    reg [7:0] z3897_assgn38970;
    reg [7:0] z3897_assgn38971;
    reg [7:0] z1351_assgn1351;
    wire [7:0]  p1ls2_G16_inv0_G256_inv0;
    wire [7:0]  e0_G256_inv0;
    wire [7:0]  e1_G256_inv0;
    wire [7:0]  r00_G16_mul1_G256_inv0;
    wire [7:0]  r10_G16_mul1_G256_inv0;
    wire [7:0]  r20_G16_mul1_G256_inv0;
    wire [7:0]  r30_G16_mul1_G256_inv0;
    wire [7:0]  r40_G16_mul1_G256_inv0;
    wire [7:0]  r50_G16_mul1_G256_inv0;
    wire [7:0]  r60_G16_mul1_G256_inv0;
    wire [7:0]  r70_G16_mul1_G256_inv0;
    wire [7:0]  r80_G16_mul1_G256_inv0;
    wire [7:0]  z3923_assgn3923;
    reg [7:0] z3923_assgn39230;
    reg [7:0] z3923_assgn39231;
    reg [7:0] z1375_assgn1375;
    wire [7:0]  a0_0_G16_mul1_G256_inv0;
    wire [7:0]  z3927_assgn3927;
    reg [7:0] z3927_assgn39270;
    reg [7:0] z3927_assgn39271;
    reg [7:0] z1377_assgn1377;
    wire [7:0]  a1_0_G16_mul1_G256_inv0;
    wire [7:0]  z3931_assgn3931;
    reg [7:0] z3931_assgn39310;
    reg [7:0] z3931_assgn39311;
    reg [7:0] z1379_assgn1379;
    wire [7:0]  a0_G16_mul1_G256_inv0;
    wire [7:0]  z3935_assgn3935;
    reg [7:0] z3935_assgn39350;
    reg [7:0] z3935_assgn39351;
    reg [7:0] z1381_assgn1381;
    wire [7:0]  a1_G16_mul1_G256_inv0;
    wire [7:0]  z3939_assgn3939;
    reg [7:0] z3939_assgn39390;
    reg [7:0] z3939_assgn39391;
    reg [7:0] z1383_assgn1383;
    wire [7:0]  b0_G16_mul1_G256_inv0;
    wire [7:0]  z3943_assgn3943;
    reg [7:0] z3943_assgn39430;
    reg [7:0] z3943_assgn39431;
    reg [7:0] z1385_assgn1385;
    wire [7:0]  b1_G16_mul1_G256_inv0;
    wire [7:0]  c0_0_G16_mul1_G256_inv0;
    wire [7:0]  c1_0_G16_mul1_G256_inv0;
    wire [7:0]  c0_G16_mul1_G256_inv0;
    wire [7:0]  c1_G16_mul1_G256_inv0;
    wire [7:0]  d0_G16_mul1_G256_inv0;
    wire [7:0]  d1_G16_mul1_G256_inv0;
    wire [7:0]  axorb_0_G16_mul1_G256_inv0;
    wire [7:0]  cxord_0_G16_mul1_G256_inv0;
    wire [7:0]  axorb_1_G16_mul1_G256_inv0;
    wire [7:0]  cxord_1_G16_mul1_G256_inv0;
    wire [7:0]  r00_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  r10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  r20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3973_assgn3973;
    reg [7:0] z3973_assgn39730;
    reg [7:0] z3973_assgn39731;
    reg [7:0] z1413_assgn1413;
    wire [7:0]  a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3977_assgn3977;
    reg [7:0] z3977_assgn39770;
    reg [7:0] z3977_assgn39771;
    reg [7:0] z1415_assgn1415;
    wire [7:0]  a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3981_assgn3981;
    reg [7:0] z3981_assgn39810;
    reg [7:0] z3981_assgn39811;
    reg [7:0] z1417_assgn1417;
    wire [7:0]  a0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3985_assgn3985;
    reg [7:0] z3985_assgn39850;
    reg [7:0] z3985_assgn39851;
    reg [7:0] z1419_assgn1419;
    wire [7:0]  a1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3989_assgn3989;
    reg [7:0] z3989_assgn39890;
    reg [7:0] z3989_assgn39891;
    reg [7:0] z1421_assgn1421;
    wire [7:0]  b0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z3993_assgn3993;
    reg [7:0] z3993_assgn39930;
    reg [7:0] z3993_assgn39931;
    reg [7:0] z1423_assgn1423;
    wire [7:0]  b1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  c0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  c1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  d0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  d1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  axorb_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4019_assgn4019;
    reg [7:0] z4019_assgn40190;
    reg [7:0] z4019_assgn40191;
    reg [7:0] z1447_assgn1447;
    wire [7:0]  p2_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4023_assgn4023;
    reg [7:0] z4023_assgn40230;
    reg [7:0] z4023_assgn40231;
    reg [7:0] z1449_assgn1449;
    wire [7:0]  i1_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4027_assgn4027;
    reg [7:0] z4027_assgn40270;
    reg [7:0] z4027_assgn40271;
    reg [7:0] z1451_assgn1451;
    wire [7:0]  p3_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4031_assgn4031;
    reg [7:0] z4031_assgn40310;
    reg [7:0] z4031_assgn40311;
    reg [7:0] z1453_assgn1453;
    wire [7:0]  i2_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4035_assgn4035;
    reg [7:0] z4035_assgn40350;
    reg [7:0] z4035_assgn40351;
    reg [7:0] z1455_assgn1455;
    wire [7:0]  p1_domand0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4039_assgn4039;
    reg [7:0] z4039_assgn40390;
    reg [7:0] z4039_assgn40391;
    reg [7:0] z1457_assgn1457;
    wire [7:0]  p4_domand0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_domand0_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  e0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_domand0_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  e1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4049_assgn4049;
    reg [7:0] z4049_assgn40490;
    reg [7:0] z4049_assgn40491;
    reg [7:0] z1465_assgn1465;
    wire [7:0]  p2_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4053_assgn4053;
    reg [7:0] z4053_assgn40530;
    reg [7:0] z4053_assgn40531;
    reg [7:0] z1467_assgn1467;
    wire [7:0]  i1_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4057_assgn4057;
    reg [7:0] z4057_assgn40570;
    reg [7:0] z4057_assgn40571;
    reg [7:0] z1469_assgn1469;
    wire [7:0]  p3_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4061_assgn4061;
    reg [7:0] z4061_assgn40610;
    reg [7:0] z4061_assgn40611;
    reg [7:0] z1471_assgn1471;
    wire [7:0]  i2_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4065_assgn4065;
    reg [7:0] z4065_assgn40650;
    reg [7:0] z4065_assgn40651;
    reg [7:0] z1473_assgn1473;
    wire [7:0]  p1_domand1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4069_assgn4069;
    reg [7:0] z4069_assgn40690;
    reg [7:0] z4069_assgn40691;
    reg [7:0] z1475_assgn1475;
    wire [7:0]  p4_domand1_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_domand1_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_domand1_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  p0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  p1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4083_assgn4083;
    reg [7:0] z4083_assgn40830;
    reg [7:0] z4083_assgn40831;
    reg [7:0] z1487_assgn1487;
    wire [7:0]  p2_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4087_assgn4087;
    reg [7:0] z4087_assgn40870;
    reg [7:0] z4087_assgn40871;
    reg [7:0] z1489_assgn1489;
    wire [7:0]  i1_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4091_assgn4091;
    reg [7:0] z4091_assgn40910;
    reg [7:0] z4091_assgn40911;
    reg [7:0] z1491_assgn1491;
    wire [7:0]  p3_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4095_assgn4095;
    reg [7:0] z4095_assgn40950;
    reg [7:0] z4095_assgn40951;
    reg [7:0] z1493_assgn1493;
    wire [7:0]  i2_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4099_assgn4099;
    reg [7:0] z4099_assgn40990;
    reg [7:0] z4099_assgn40991;
    reg [7:0] z1495_assgn1495;
    wire [7:0]  p1_domand2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4103_assgn4103;
    reg [7:0] z4103_assgn41030;
    reg [7:0] z4103_assgn41031;
    reg [7:0] z1497_assgn1497;
    wire [7:0]  p4_domand2_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i1_domand2_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] i2_domand2_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  q0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  q1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4115_assgn4115;
    reg [7:0] z4115_assgn41150;
    reg [7:0] z4115_assgn41151;
    reg [7:0] z4115_assgn41152;
    reg [7:0] z1507_assgn1507;
    wire [7:0]  p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  z4119_assgn4119;
    reg [7:0] z4119_assgn41190;
    reg [7:0] z4119_assgn41191;
    reg [7:0] z4119_assgn41192;
    reg [7:0] z1509_assgn1509;
    wire [7:0]  p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0]  e0_G16_mul1_G256_inv0;
    wire [7:0]  e1_G16_mul1_G256_inv0;
    wire [7:0]  z4127_assgn4127;
    reg [7:0] z4127_assgn41270;
    reg [7:0] z4127_assgn41271;
    reg [7:0] z4127_assgn41272;
    reg [7:0] z1515_assgn1515;
    wire [7:0]  a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4131_assgn4131;
    reg [7:0] z4131_assgn41310;
    reg [7:0] z4131_assgn41311;
    reg [7:0] z4131_assgn41312;
    reg [7:0] z1517_assgn1517;
    wire [7:0]  a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4135_assgn4135;
    reg [7:0] z4135_assgn41350;
    reg [7:0] z4135_assgn41351;
    reg [7:0] z4135_assgn41352;
    reg [7:0] z1519_assgn1519;
    wire [7:0]  a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4139_assgn4139;
    reg [7:0] z4139_assgn41390;
    reg [7:0] z4139_assgn41391;
    reg [7:0] z4139_assgn41392;
    reg [7:0] z1521_assgn1521;
    wire [7:0]  a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4143_assgn4143;
    reg [7:0] z4143_assgn41430;
    reg [7:0] z4143_assgn41431;
    reg [7:0] z4143_assgn41432;
    reg [7:0] z1523_assgn1523;
    wire [7:0]  b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4147_assgn4147;
    reg [7:0] z4147_assgn41470;
    reg [7:0] z4147_assgn41471;
    reg [7:0] z4147_assgn41472;
    reg [7:0] z1525_assgn1525;
    wire [7:0]  b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4159_assgn4159;
    reg [7:0] z4159_assgn41590;
    reg [7:0] z4159_assgn41591;
    reg [7:0] z4159_assgn41592;
    reg [7:0] z1535_assgn1535;
    wire [7:0]  p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  z4163_assgn4163;
    reg [7:0] z4163_assgn41630;
    reg [7:0] z4163_assgn41631;
    reg [7:0] z4163_assgn41632;
    reg [7:0] z1537_assgn1537;
    wire [7:0]  p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0]  e01_G16_mul1_G256_inv0;
    wire [7:0]  e11_G16_mul1_G256_inv0;
    wire [7:0]  r00_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  r10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  r20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4177_assgn4177;
    reg [7:0] z4177_assgn41770;
    reg [7:0] z4177_assgn41771;
    reg [7:0] z1549_assgn1549;
    wire [7:0]  a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4181_assgn4181;
    reg [7:0] z4181_assgn41810;
    reg [7:0] z4181_assgn41811;
    reg [7:0] z1551_assgn1551;
    wire [7:0]  a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4185_assgn4185;
    reg [7:0] z4185_assgn41850;
    reg [7:0] z4185_assgn41851;
    reg [7:0] z1553_assgn1553;
    wire [7:0]  a0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4189_assgn4189;
    reg [7:0] z4189_assgn41890;
    reg [7:0] z4189_assgn41891;
    reg [7:0] z1555_assgn1555;
    wire [7:0]  a1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4193_assgn4193;
    reg [7:0] z4193_assgn41930;
    reg [7:0] z4193_assgn41931;
    reg [7:0] z1557_assgn1557;
    wire [7:0]  b0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4197_assgn4197;
    reg [7:0] z4197_assgn41970;
    reg [7:0] z4197_assgn41971;
    reg [7:0] z1559_assgn1559;
    wire [7:0]  b1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  c0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  c1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  d0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  d1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  axorb_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4223_assgn4223;
    reg [7:0] z4223_assgn42230;
    reg [7:0] z4223_assgn42231;
    reg [7:0] z1583_assgn1583;
    wire [7:0]  p2_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4227_assgn4227;
    reg [7:0] z4227_assgn42270;
    reg [7:0] z4227_assgn42271;
    reg [7:0] z1585_assgn1585;
    wire [7:0]  i1_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4231_assgn4231;
    reg [7:0] z4231_assgn42310;
    reg [7:0] z4231_assgn42311;
    reg [7:0] z1587_assgn1587;
    wire [7:0]  p3_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4235_assgn4235;
    reg [7:0] z4235_assgn42350;
    reg [7:0] z4235_assgn42351;
    reg [7:0] z1589_assgn1589;
    wire [7:0]  i2_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4239_assgn4239;
    reg [7:0] z4239_assgn42390;
    reg [7:0] z4239_assgn42391;
    reg [7:0] z1591_assgn1591;
    wire [7:0]  p1_domand0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4243_assgn4243;
    reg [7:0] z4243_assgn42430;
    reg [7:0] z4243_assgn42431;
    reg [7:0] z1593_assgn1593;
    wire [7:0]  p4_domand0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_domand0_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  e0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_domand0_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  e1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4253_assgn4253;
    reg [7:0] z4253_assgn42530;
    reg [7:0] z4253_assgn42531;
    reg [7:0] z1601_assgn1601;
    wire [7:0]  p2_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4257_assgn4257;
    reg [7:0] z4257_assgn42570;
    reg [7:0] z4257_assgn42571;
    reg [7:0] z1603_assgn1603;
    wire [7:0]  i1_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4261_assgn4261;
    reg [7:0] z4261_assgn42610;
    reg [7:0] z4261_assgn42611;
    reg [7:0] z1605_assgn1605;
    wire [7:0]  p3_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4265_assgn4265;
    reg [7:0] z4265_assgn42650;
    reg [7:0] z4265_assgn42651;
    reg [7:0] z1607_assgn1607;
    wire [7:0]  i2_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4269_assgn4269;
    reg [7:0] z4269_assgn42690;
    reg [7:0] z4269_assgn42691;
    reg [7:0] z1609_assgn1609;
    wire [7:0]  p1_domand1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4273_assgn4273;
    reg [7:0] z4273_assgn42730;
    reg [7:0] z4273_assgn42731;
    reg [7:0] z1611_assgn1611;
    wire [7:0]  p4_domand1_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_domand1_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_domand1_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  p0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  p1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4287_assgn4287;
    reg [7:0] z4287_assgn42870;
    reg [7:0] z4287_assgn42871;
    reg [7:0] z1623_assgn1623;
    wire [7:0]  p2_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4291_assgn4291;
    reg [7:0] z4291_assgn42910;
    reg [7:0] z4291_assgn42911;
    reg [7:0] z1625_assgn1625;
    wire [7:0]  i1_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4295_assgn4295;
    reg [7:0] z4295_assgn42950;
    reg [7:0] z4295_assgn42951;
    reg [7:0] z1627_assgn1627;
    wire [7:0]  p3_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4299_assgn4299;
    reg [7:0] z4299_assgn42990;
    reg [7:0] z4299_assgn42991;
    reg [7:0] z1629_assgn1629;
    wire [7:0]  i2_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4303_assgn4303;
    reg [7:0] z4303_assgn43030;
    reg [7:0] z4303_assgn43031;
    reg [7:0] z1631_assgn1631;
    wire [7:0]  p1_domand2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4307_assgn4307;
    reg [7:0] z4307_assgn43070;
    reg [7:0] z4307_assgn43071;
    reg [7:0] z1633_assgn1633;
    wire [7:0]  p4_domand2_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i1_domand2_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] i2_domand2_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  q0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  q1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4319_assgn4319;
    reg [7:0] z4319_assgn43190;
    reg [7:0] z4319_assgn43191;
    reg [7:0] z4319_assgn43192;
    reg [7:0] z1643_assgn1643;
    wire [7:0]  p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  z4323_assgn4323;
    reg [7:0] z4323_assgn43230;
    reg [7:0] z4323_assgn43231;
    reg [7:0] z4323_assgn43232;
    reg [7:0] z1645_assgn1645;
    wire [7:0]  p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0]  p0_0_G16_mul1_G256_inv0;
    wire [7:0]  p1_0_G16_mul1_G256_inv0;
    wire [7:0]  p0_G16_mul1_G256_inv0;
    wire [7:0]  p1_G16_mul1_G256_inv0;
    wire [7:0]  r00_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  r10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  r20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4341_assgn4341;
    reg [7:0] z4341_assgn43410;
    reg [7:0] z4341_assgn43411;
    reg [7:0] z1661_assgn1661;
    wire [7:0]  a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4345_assgn4345;
    reg [7:0] z4345_assgn43450;
    reg [7:0] z4345_assgn43451;
    reg [7:0] z1663_assgn1663;
    wire [7:0]  a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4349_assgn4349;
    reg [7:0] z4349_assgn43490;
    reg [7:0] z4349_assgn43491;
    reg [7:0] z1665_assgn1665;
    wire [7:0]  a0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4353_assgn4353;
    reg [7:0] z4353_assgn43530;
    reg [7:0] z4353_assgn43531;
    reg [7:0] z1667_assgn1667;
    wire [7:0]  a1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4357_assgn4357;
    reg [7:0] z4357_assgn43570;
    reg [7:0] z4357_assgn43571;
    reg [7:0] z1669_assgn1669;
    wire [7:0]  b0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4361_assgn4361;
    reg [7:0] z4361_assgn43610;
    reg [7:0] z4361_assgn43611;
    reg [7:0] z1671_assgn1671;
    wire [7:0]  b1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  c0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  c1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  d0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  d1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  axorb_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4387_assgn4387;
    reg [7:0] z4387_assgn43870;
    reg [7:0] z4387_assgn43871;
    reg [7:0] z1695_assgn1695;
    wire [7:0]  p2_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4391_assgn4391;
    reg [7:0] z4391_assgn43910;
    reg [7:0] z4391_assgn43911;
    reg [7:0] z1697_assgn1697;
    wire [7:0]  i1_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4395_assgn4395;
    reg [7:0] z4395_assgn43950;
    reg [7:0] z4395_assgn43951;
    reg [7:0] z1699_assgn1699;
    wire [7:0]  p3_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4399_assgn4399;
    reg [7:0] z4399_assgn43990;
    reg [7:0] z4399_assgn43991;
    reg [7:0] z1701_assgn1701;
    wire [7:0]  i2_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4403_assgn4403;
    reg [7:0] z4403_assgn44030;
    reg [7:0] z4403_assgn44031;
    reg [7:0] z1703_assgn1703;
    wire [7:0]  p1_domand0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4407_assgn4407;
    reg [7:0] z4407_assgn44070;
    reg [7:0] z4407_assgn44071;
    reg [7:0] z1705_assgn1705;
    wire [7:0]  p4_domand0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_domand0_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  e0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_domand0_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  e1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4417_assgn4417;
    reg [7:0] z4417_assgn44170;
    reg [7:0] z4417_assgn44171;
    reg [7:0] z1713_assgn1713;
    wire [7:0]  p2_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4421_assgn4421;
    reg [7:0] z4421_assgn44210;
    reg [7:0] z4421_assgn44211;
    reg [7:0] z1715_assgn1715;
    wire [7:0]  i1_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4425_assgn4425;
    reg [7:0] z4425_assgn44250;
    reg [7:0] z4425_assgn44251;
    reg [7:0] z1717_assgn1717;
    wire [7:0]  p3_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4429_assgn4429;
    reg [7:0] z4429_assgn44290;
    reg [7:0] z4429_assgn44291;
    reg [7:0] z1719_assgn1719;
    wire [7:0]  i2_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4433_assgn4433;
    reg [7:0] z4433_assgn44330;
    reg [7:0] z4433_assgn44331;
    reg [7:0] z1721_assgn1721;
    wire [7:0]  p1_domand1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4437_assgn4437;
    reg [7:0] z4437_assgn44370;
    reg [7:0] z4437_assgn44371;
    reg [7:0] z1723_assgn1723;
    wire [7:0]  p4_domand1_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_domand1_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_domand1_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  p0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  p1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4451_assgn4451;
    reg [7:0] z4451_assgn44510;
    reg [7:0] z4451_assgn44511;
    reg [7:0] z1735_assgn1735;
    wire [7:0]  p2_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4455_assgn4455;
    reg [7:0] z4455_assgn44550;
    reg [7:0] z4455_assgn44551;
    reg [7:0] z1737_assgn1737;
    wire [7:0]  i1_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4459_assgn4459;
    reg [7:0] z4459_assgn44590;
    reg [7:0] z4459_assgn44591;
    reg [7:0] z1739_assgn1739;
    wire [7:0]  p3_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4463_assgn4463;
    reg [7:0] z4463_assgn44630;
    reg [7:0] z4463_assgn44631;
    reg [7:0] z1741_assgn1741;
    wire [7:0]  i2_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4467_assgn4467;
    reg [7:0] z4467_assgn44670;
    reg [7:0] z4467_assgn44671;
    reg [7:0] z1743_assgn1743;
    wire [7:0]  p1_domand2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4471_assgn4471;
    reg [7:0] z4471_assgn44710;
    reg [7:0] z4471_assgn44711;
    reg [7:0] z1745_assgn1745;
    wire [7:0]  p4_domand2_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i1_domand2_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] i2_domand2_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  q0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  q1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4483_assgn4483;
    reg [7:0] z4483_assgn44830;
    reg [7:0] z4483_assgn44831;
    reg [7:0] z4483_assgn44832;
    reg [7:0] z1755_assgn1755;
    wire [7:0]  p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  z4487_assgn4487;
    reg [7:0] z4487_assgn44870;
    reg [7:0] z4487_assgn44871;
    reg [7:0] z4487_assgn44872;
    reg [7:0] z1757_assgn1757;
    wire [7:0]  p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0]  q0_0_G16_mul1_G256_inv0;
    wire [7:0]  q1_0_G16_mul1_G256_inv0;
    wire [7:0]  q0_G16_mul1_G256_inv0;
    wire [7:0]  q1_G16_mul1_G256_inv0;
    wire [7:0]  z4499_assgn4499;
    reg [7:0] z4499_assgn44990;
    reg [7:0] z4499_assgn44991;
    reg [7:0] z4499_assgn44992;
    reg [7:0] z1767_assgn1767;
    wire [7:0]  p0ls2_G16_mul1_G256_inv0;
    wire [7:0]  z4503_assgn4503;
    reg [7:0] z4503_assgn45030;
    reg [7:0] z4503_assgn45031;
    reg [7:0] z4503_assgn45032;
    reg [7:0] z1769_assgn1769;
    wire [7:0]  p1ls2_G16_mul1_G256_inv0;
    wire [7:0]  p0_G256_inv0;
    wire [7:0]  p1_G256_inv0;
    wire [7:0]  r00_G16_mul2_G256_inv0;
    wire [7:0]  r10_G16_mul2_G256_inv0;
    wire [7:0]  r20_G16_mul2_G256_inv0;
    wire [7:0]  r30_G16_mul2_G256_inv0;
    wire [7:0]  r40_G16_mul2_G256_inv0;
    wire [7:0]  r50_G16_mul2_G256_inv0;
    wire [7:0]  r60_G16_mul2_G256_inv0;
    wire [7:0]  r70_G16_mul2_G256_inv0;
    wire [7:0]  r80_G16_mul2_G256_inv0;
    wire [7:0]  z4529_assgn4529;
    reg [7:0] z4529_assgn45290;
    reg [7:0] z4529_assgn45291;
    reg [7:0] z1793_assgn1793;
    wire [7:0]  a0_0_G16_mul2_G256_inv0;
    wire [7:0]  z4533_assgn4533;
    reg [7:0] z4533_assgn45330;
    reg [7:0] z4533_assgn45331;
    reg [7:0] z1795_assgn1795;
    wire [7:0]  a1_0_G16_mul2_G256_inv0;
    wire [7:0]  z4537_assgn4537;
    reg [7:0] z4537_assgn45370;
    reg [7:0] z4537_assgn45371;
    reg [7:0] z1797_assgn1797;
    wire [7:0]  a0_G16_mul2_G256_inv0;
    wire [7:0]  z4541_assgn4541;
    reg [7:0] z4541_assgn45410;
    reg [7:0] z4541_assgn45411;
    reg [7:0] z1799_assgn1799;
    wire [7:0]  a1_G16_mul2_G256_inv0;
    wire [7:0]  z4545_assgn4545;
    reg [7:0] z4545_assgn45450;
    reg [7:0] z4545_assgn45451;
    reg [7:0] z1801_assgn1801;
    wire [7:0]  b0_G16_mul2_G256_inv0;
    wire [7:0]  z4549_assgn4549;
    reg [7:0] z4549_assgn45490;
    reg [7:0] z4549_assgn45491;
    reg [7:0] z1803_assgn1803;
    wire [7:0]  b1_G16_mul2_G256_inv0;
    wire [7:0]  c0_0_G16_mul2_G256_inv0;
    wire [7:0]  c1_0_G16_mul2_G256_inv0;
    wire [7:0]  c0_G16_mul2_G256_inv0;
    wire [7:0]  c1_G16_mul2_G256_inv0;
    wire [7:0]  d0_G16_mul2_G256_inv0;
    wire [7:0]  d1_G16_mul2_G256_inv0;
    wire [7:0]  axorb_0_G16_mul2_G256_inv0;
    wire [7:0]  cxord_0_G16_mul2_G256_inv0;
    wire [7:0]  axorb_1_G16_mul2_G256_inv0;
    wire [7:0]  cxord_1_G16_mul2_G256_inv0;
    wire [7:0]  r00_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  r10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  r20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4579_assgn4579;
    reg [7:0] z4579_assgn45790;
    reg [7:0] z4579_assgn45791;
    reg [7:0] z1831_assgn1831;
    wire [7:0]  a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4583_assgn4583;
    reg [7:0] z4583_assgn45830;
    reg [7:0] z4583_assgn45831;
    reg [7:0] z1833_assgn1833;
    wire [7:0]  a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4587_assgn4587;
    reg [7:0] z4587_assgn45870;
    reg [7:0] z4587_assgn45871;
    reg [7:0] z1835_assgn1835;
    wire [7:0]  a0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4591_assgn4591;
    reg [7:0] z4591_assgn45910;
    reg [7:0] z4591_assgn45911;
    reg [7:0] z1837_assgn1837;
    wire [7:0]  a1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4595_assgn4595;
    reg [7:0] z4595_assgn45950;
    reg [7:0] z4595_assgn45951;
    reg [7:0] z1839_assgn1839;
    wire [7:0]  b0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4599_assgn4599;
    reg [7:0] z4599_assgn45990;
    reg [7:0] z4599_assgn45991;
    reg [7:0] z1841_assgn1841;
    wire [7:0]  b1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  c0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  c1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  d0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  d1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  axorb_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4625_assgn4625;
    reg [7:0] z4625_assgn46250;
    reg [7:0] z4625_assgn46251;
    reg [7:0] z1865_assgn1865;
    wire [7:0]  p2_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4629_assgn4629;
    reg [7:0] z4629_assgn46290;
    reg [7:0] z4629_assgn46291;
    reg [7:0] z1867_assgn1867;
    wire [7:0]  i1_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4633_assgn4633;
    reg [7:0] z4633_assgn46330;
    reg [7:0] z4633_assgn46331;
    reg [7:0] z1869_assgn1869;
    wire [7:0]  p3_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4637_assgn4637;
    reg [7:0] z4637_assgn46370;
    reg [7:0] z4637_assgn46371;
    reg [7:0] z1871_assgn1871;
    wire [7:0]  i2_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4641_assgn4641;
    reg [7:0] z4641_assgn46410;
    reg [7:0] z4641_assgn46411;
    reg [7:0] z1873_assgn1873;
    wire [7:0]  p1_domand0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4645_assgn4645;
    reg [7:0] z4645_assgn46450;
    reg [7:0] z4645_assgn46451;
    reg [7:0] z1875_assgn1875;
    wire [7:0]  p4_domand0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_domand0_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  e0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_domand0_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  e1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4655_assgn4655;
    reg [7:0] z4655_assgn46550;
    reg [7:0] z4655_assgn46551;
    reg [7:0] z1883_assgn1883;
    wire [7:0]  p2_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4659_assgn4659;
    reg [7:0] z4659_assgn46590;
    reg [7:0] z4659_assgn46591;
    reg [7:0] z1885_assgn1885;
    wire [7:0]  i1_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4663_assgn4663;
    reg [7:0] z4663_assgn46630;
    reg [7:0] z4663_assgn46631;
    reg [7:0] z1887_assgn1887;
    wire [7:0]  p3_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4667_assgn4667;
    reg [7:0] z4667_assgn46670;
    reg [7:0] z4667_assgn46671;
    reg [7:0] z1889_assgn1889;
    wire [7:0]  i2_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4671_assgn4671;
    reg [7:0] z4671_assgn46710;
    reg [7:0] z4671_assgn46711;
    reg [7:0] z1891_assgn1891;
    wire [7:0]  p1_domand1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4675_assgn4675;
    reg [7:0] z4675_assgn46750;
    reg [7:0] z4675_assgn46751;
    reg [7:0] z1893_assgn1893;
    wire [7:0]  p4_domand1_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_domand1_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_domand1_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  p0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  p1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4689_assgn4689;
    reg [7:0] z4689_assgn46890;
    reg [7:0] z4689_assgn46891;
    reg [7:0] z1905_assgn1905;
    wire [7:0]  p2_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4693_assgn4693;
    reg [7:0] z4693_assgn46930;
    reg [7:0] z4693_assgn46931;
    reg [7:0] z1907_assgn1907;
    wire [7:0]  i1_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4697_assgn4697;
    reg [7:0] z4697_assgn46970;
    reg [7:0] z4697_assgn46971;
    reg [7:0] z1909_assgn1909;
    wire [7:0]  p3_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4701_assgn4701;
    reg [7:0] z4701_assgn47010;
    reg [7:0] z4701_assgn47011;
    reg [7:0] z1911_assgn1911;
    wire [7:0]  i2_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4705_assgn4705;
    reg [7:0] z4705_assgn47050;
    reg [7:0] z4705_assgn47051;
    reg [7:0] z1913_assgn1913;
    wire [7:0]  p1_domand2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4709_assgn4709;
    reg [7:0] z4709_assgn47090;
    reg [7:0] z4709_assgn47091;
    reg [7:0] z1915_assgn1915;
    wire [7:0]  p4_domand2_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i1_domand2_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] i2_domand2_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  q0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  q1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4721_assgn4721;
    reg [7:0] z4721_assgn47210;
    reg [7:0] z4721_assgn47211;
    reg [7:0] z4721_assgn47212;
    reg [7:0] z1925_assgn1925;
    wire [7:0]  p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  z4725_assgn4725;
    reg [7:0] z4725_assgn47250;
    reg [7:0] z4725_assgn47251;
    reg [7:0] z4725_assgn47252;
    reg [7:0] z1927_assgn1927;
    wire [7:0]  p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0]  e0_G16_mul2_G256_inv0;
    wire [7:0]  e1_G16_mul2_G256_inv0;
    wire [7:0]  z4733_assgn4733;
    reg [7:0] z4733_assgn47330;
    reg [7:0] z4733_assgn47331;
    reg [7:0] z4733_assgn47332;
    reg [7:0] z1933_assgn1933;
    wire [7:0]  a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4737_assgn4737;
    reg [7:0] z4737_assgn47370;
    reg [7:0] z4737_assgn47371;
    reg [7:0] z4737_assgn47372;
    reg [7:0] z1935_assgn1935;
    wire [7:0]  a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4741_assgn4741;
    reg [7:0] z4741_assgn47410;
    reg [7:0] z4741_assgn47411;
    reg [7:0] z4741_assgn47412;
    reg [7:0] z1937_assgn1937;
    wire [7:0]  a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4745_assgn4745;
    reg [7:0] z4745_assgn47450;
    reg [7:0] z4745_assgn47451;
    reg [7:0] z4745_assgn47452;
    reg [7:0] z1939_assgn1939;
    wire [7:0]  a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4749_assgn4749;
    reg [7:0] z4749_assgn47490;
    reg [7:0] z4749_assgn47491;
    reg [7:0] z4749_assgn47492;
    reg [7:0] z1941_assgn1941;
    wire [7:0]  b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4753_assgn4753;
    reg [7:0] z4753_assgn47530;
    reg [7:0] z4753_assgn47531;
    reg [7:0] z4753_assgn47532;
    reg [7:0] z1943_assgn1943;
    wire [7:0]  b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4765_assgn4765;
    reg [7:0] z4765_assgn47650;
    reg [7:0] z4765_assgn47651;
    reg [7:0] z4765_assgn47652;
    reg [7:0] z1953_assgn1953;
    wire [7:0]  p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  z4769_assgn4769;
    reg [7:0] z4769_assgn47690;
    reg [7:0] z4769_assgn47691;
    reg [7:0] z4769_assgn47692;
    reg [7:0] z1955_assgn1955;
    wire [7:0]  p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0]  e01_G16_mul2_G256_inv0;
    wire [7:0]  e11_G16_mul2_G256_inv0;
    wire [7:0]  r00_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  r10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  r20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4783_assgn4783;
    reg [7:0] z4783_assgn47830;
    reg [7:0] z4783_assgn47831;
    reg [7:0] z1967_assgn1967;
    wire [7:0]  a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4787_assgn4787;
    reg [7:0] z4787_assgn47870;
    reg [7:0] z4787_assgn47871;
    reg [7:0] z1969_assgn1969;
    wire [7:0]  a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4791_assgn4791;
    reg [7:0] z4791_assgn47910;
    reg [7:0] z4791_assgn47911;
    reg [7:0] z1971_assgn1971;
    wire [7:0]  a0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4795_assgn4795;
    reg [7:0] z4795_assgn47950;
    reg [7:0] z4795_assgn47951;
    reg [7:0] z1973_assgn1973;
    wire [7:0]  a1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4799_assgn4799;
    reg [7:0] z4799_assgn47990;
    reg [7:0] z4799_assgn47991;
    reg [7:0] z1975_assgn1975;
    wire [7:0]  b0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4803_assgn4803;
    reg [7:0] z4803_assgn48030;
    reg [7:0] z4803_assgn48031;
    reg [7:0] z1977_assgn1977;
    wire [7:0]  b1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  c0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  c1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  d0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  d1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  axorb_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4829_assgn4829;
    reg [7:0] z4829_assgn48290;
    reg [7:0] z4829_assgn48291;
    reg [7:0] z2001_assgn2001;
    wire [7:0]  p2_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4833_assgn4833;
    reg [7:0] z4833_assgn48330;
    reg [7:0] z4833_assgn48331;
    reg [7:0] z2003_assgn2003;
    wire [7:0]  i1_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4837_assgn4837;
    reg [7:0] z4837_assgn48370;
    reg [7:0] z4837_assgn48371;
    reg [7:0] z2005_assgn2005;
    wire [7:0]  p3_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4841_assgn4841;
    reg [7:0] z4841_assgn48410;
    reg [7:0] z4841_assgn48411;
    reg [7:0] z2007_assgn2007;
    wire [7:0]  i2_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4845_assgn4845;
    reg [7:0] z4845_assgn48450;
    reg [7:0] z4845_assgn48451;
    reg [7:0] z2009_assgn2009;
    wire [7:0]  p1_domand0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4849_assgn4849;
    reg [7:0] z4849_assgn48490;
    reg [7:0] z4849_assgn48491;
    reg [7:0] z2011_assgn2011;
    wire [7:0]  p4_domand0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_domand0_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  e0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_domand0_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  e1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4859_assgn4859;
    reg [7:0] z4859_assgn48590;
    reg [7:0] z4859_assgn48591;
    reg [7:0] z2019_assgn2019;
    wire [7:0]  p2_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4863_assgn4863;
    reg [7:0] z4863_assgn48630;
    reg [7:0] z4863_assgn48631;
    reg [7:0] z2021_assgn2021;
    wire [7:0]  i1_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4867_assgn4867;
    reg [7:0] z4867_assgn48670;
    reg [7:0] z4867_assgn48671;
    reg [7:0] z2023_assgn2023;
    wire [7:0]  p3_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4871_assgn4871;
    reg [7:0] z4871_assgn48710;
    reg [7:0] z4871_assgn48711;
    reg [7:0] z2025_assgn2025;
    wire [7:0]  i2_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4875_assgn4875;
    reg [7:0] z4875_assgn48750;
    reg [7:0] z4875_assgn48751;
    reg [7:0] z2027_assgn2027;
    wire [7:0]  p1_domand1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4879_assgn4879;
    reg [7:0] z4879_assgn48790;
    reg [7:0] z4879_assgn48791;
    reg [7:0] z2029_assgn2029;
    wire [7:0]  p4_domand1_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_domand1_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_domand1_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  p0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  p1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4893_assgn4893;
    reg [7:0] z4893_assgn48930;
    reg [7:0] z4893_assgn48931;
    reg [7:0] z2041_assgn2041;
    wire [7:0]  p2_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4897_assgn4897;
    reg [7:0] z4897_assgn48970;
    reg [7:0] z4897_assgn48971;
    reg [7:0] z2043_assgn2043;
    wire [7:0]  i1_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4901_assgn4901;
    reg [7:0] z4901_assgn49010;
    reg [7:0] z4901_assgn49011;
    reg [7:0] z2045_assgn2045;
    wire [7:0]  p3_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4905_assgn4905;
    reg [7:0] z4905_assgn49050;
    reg [7:0] z4905_assgn49051;
    reg [7:0] z2047_assgn2047;
    wire [7:0]  i2_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4909_assgn4909;
    reg [7:0] z4909_assgn49090;
    reg [7:0] z4909_assgn49091;
    reg [7:0] z2049_assgn2049;
    wire [7:0]  p1_domand2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4913_assgn4913;
    reg [7:0] z4913_assgn49130;
    reg [7:0] z4913_assgn49131;
    reg [7:0] z2051_assgn2051;
    wire [7:0]  p4_domand2_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i1_domand2_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] i2_domand2_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  q0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  q1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4925_assgn4925;
    reg [7:0] z4925_assgn49250;
    reg [7:0] z4925_assgn49251;
    reg [7:0] z4925_assgn49252;
    reg [7:0] z2061_assgn2061;
    wire [7:0]  p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  z4929_assgn4929;
    reg [7:0] z4929_assgn49290;
    reg [7:0] z4929_assgn49291;
    reg [7:0] z4929_assgn49292;
    reg [7:0] z2063_assgn2063;
    wire [7:0]  p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0]  p0_0_G16_mul2_G256_inv0;
    wire [7:0]  p1_0_G16_mul2_G256_inv0;
    wire [7:0]  p0_G16_mul2_G256_inv0;
    wire [7:0]  p1_G16_mul2_G256_inv0;
    wire [7:0]  r00_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  r10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  r20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4947_assgn4947;
    reg [7:0] z4947_assgn49470;
    reg [7:0] z4947_assgn49471;
    reg [7:0] z2079_assgn2079;
    wire [7:0]  a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4951_assgn4951;
    reg [7:0] z4951_assgn49510;
    reg [7:0] z4951_assgn49511;
    reg [7:0] z2081_assgn2081;
    wire [7:0]  a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4955_assgn4955;
    reg [7:0] z4955_assgn49550;
    reg [7:0] z4955_assgn49551;
    reg [7:0] z2083_assgn2083;
    wire [7:0]  a0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4959_assgn4959;
    reg [7:0] z4959_assgn49590;
    reg [7:0] z4959_assgn49591;
    reg [7:0] z2085_assgn2085;
    wire [7:0]  a1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4963_assgn4963;
    reg [7:0] z4963_assgn49630;
    reg [7:0] z4963_assgn49631;
    reg [7:0] z2087_assgn2087;
    wire [7:0]  b0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4967_assgn4967;
    reg [7:0] z4967_assgn49670;
    reg [7:0] z4967_assgn49671;
    reg [7:0] z2089_assgn2089;
    wire [7:0]  b1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  c0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  c1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  d0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  d1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  axorb_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4993_assgn4993;
    reg [7:0] z4993_assgn49930;
    reg [7:0] z4993_assgn49931;
    reg [7:0] z2113_assgn2113;
    wire [7:0]  p2_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z4997_assgn4997;
    reg [7:0] z4997_assgn49970;
    reg [7:0] z4997_assgn49971;
    reg [7:0] z2115_assgn2115;
    wire [7:0]  i1_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5001_assgn5001;
    reg [7:0] z5001_assgn50010;
    reg [7:0] z5001_assgn50011;
    reg [7:0] z2117_assgn2117;
    wire [7:0]  p3_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5005_assgn5005;
    reg [7:0] z5005_assgn50050;
    reg [7:0] z5005_assgn50051;
    reg [7:0] z2119_assgn2119;
    wire [7:0]  i2_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5009_assgn5009;
    reg [7:0] z5009_assgn50090;
    reg [7:0] z5009_assgn50091;
    reg [7:0] z2121_assgn2121;
    wire [7:0]  p1_domand0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5013_assgn5013;
    reg [7:0] z5013_assgn50130;
    reg [7:0] z5013_assgn50131;
    reg [7:0] z2123_assgn2123;
    wire [7:0]  p4_domand0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_domand0_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  e0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_domand0_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  e1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5023_assgn5023;
    reg [7:0] z5023_assgn50230;
    reg [7:0] z5023_assgn50231;
    reg [7:0] z2131_assgn2131;
    wire [7:0]  p2_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5027_assgn5027;
    reg [7:0] z5027_assgn50270;
    reg [7:0] z5027_assgn50271;
    reg [7:0] z2133_assgn2133;
    wire [7:0]  i1_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5031_assgn5031;
    reg [7:0] z5031_assgn50310;
    reg [7:0] z5031_assgn50311;
    reg [7:0] z2135_assgn2135;
    wire [7:0]  p3_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5035_assgn5035;
    reg [7:0] z5035_assgn50350;
    reg [7:0] z5035_assgn50351;
    reg [7:0] z2137_assgn2137;
    wire [7:0]  i2_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5039_assgn5039;
    reg [7:0] z5039_assgn50390;
    reg [7:0] z5039_assgn50391;
    reg [7:0] z2139_assgn2139;
    wire [7:0]  p1_domand1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5043_assgn5043;
    reg [7:0] z5043_assgn50430;
    reg [7:0] z5043_assgn50431;
    reg [7:0] z2141_assgn2141;
    wire [7:0]  p4_domand1_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_domand1_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  p0_0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_domand1_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  p0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  p1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z0_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5057_assgn5057;
    reg [7:0] z5057_assgn50570;
    reg [7:0] z5057_assgn50571;
    reg [7:0] z2153_assgn2153;
    wire [7:0]  p2_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5061_assgn5061;
    reg [7:0] z5061_assgn50610;
    reg [7:0] z5061_assgn50611;
    reg [7:0] z2155_assgn2155;
    wire [7:0]  i1_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5065_assgn5065;
    reg [7:0] z5065_assgn50650;
    reg [7:0] z5065_assgn50651;
    reg [7:0] z2157_assgn2157;
    wire [7:0]  p3_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5069_assgn5069;
    reg [7:0] z5069_assgn50690;
    reg [7:0] z5069_assgn50691;
    reg [7:0] z2159_assgn2159;
    wire [7:0]  i2_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5073_assgn5073;
    reg [7:0] z5073_assgn50730;
    reg [7:0] z5073_assgn50731;
    reg [7:0] z2161_assgn2161;
    wire [7:0]  p1_domand2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5077_assgn5077;
    reg [7:0] z5077_assgn50770;
    reg [7:0] z5077_assgn50771;
    reg [7:0] z2163_assgn2163;
    wire [7:0]  p4_domand2_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i1_domand2_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_domand2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  q0_0_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] i2_domand2_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p4_domand2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0]  q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  q0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  q1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5089_assgn5089;
    reg [7:0] z5089_assgn50890;
    reg [7:0] z5089_assgn50891;
    reg [7:0] z5089_assgn50892;
    reg [7:0] z2173_assgn2173;
    wire [7:0]  p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  z5093_assgn5093;
    reg [7:0] z5093_assgn50930;
    reg [7:0] z5093_assgn50931;
    reg [7:0] z5093_assgn50932;
    reg [7:0] z2175_assgn2175;
    wire [7:0]  p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0]  q0_0_G16_mul2_G256_inv0;
    wire [7:0]  q1_0_G16_mul2_G256_inv0;
    wire [7:0]  q0_G16_mul2_G256_inv0;
    wire [7:0]  q1_G16_mul2_G256_inv0;
    wire [7:0]  z5105_assgn5105;
    reg [7:0] z5105_assgn51050;
    reg [7:0] z5105_assgn51051;
    reg [7:0] z5105_assgn51052;
    reg [7:0] z2185_assgn2185;
    wire [7:0]  p0ls2_G16_mul2_G256_inv0;
    wire [7:0]  z5109_assgn5109;
    reg [7:0] z5109_assgn51090;
    reg [7:0] z5109_assgn51091;
    reg [7:0] z5109_assgn51092;
    reg [7:0] z2187_assgn2187;
    wire [7:0]  p1ls2_G16_mul2_G256_inv0;
    wire [7:0]  q0_G256_inv0;
    wire [7:0]  q1_G256_inv0;
    wire [7:0]  z5117_assgn5117;
    reg [7:0] z5117_assgn51170;
    reg [7:0] z5117_assgn51171;
    reg [7:0] z5117_assgn51172;
    reg [7:0] z2193_assgn2193;
    wire [7:0]  p0ls4_G256_inv0;
    wire [7:0]  z5121_assgn5121;
    reg [7:0] z5121_assgn51210;
    reg [7:0] z5121_assgn51211;
    reg [7:0] z5121_assgn51212;
    reg [7:0] z2195_assgn2195;
    wire [7:0]  p1ls4_G256_inv0;
    wire [7:0]  t4;
    wire [7:0]  t5;
    wire [7:0]  y_G256_newbasis1;
    wire [7:0]  tempy1_G256_newbasis1;
    wire [7:0]  z5133_assgn5133;
    reg [7:0] z5133_assgn51330;
    reg [7:0] z5133_assgn51331;
    reg [7:0] z5133_assgn51332;
    reg [7:0] z2205_assgn2205;
    wire [7:0]  cond1_G256_newbasis1;
    wire [7:0]  negCond1_G256_newbasis1;
    wire [7:0]  yxorb1_G256_newbasis1;
    wire [7:0]  z5141_assgn5141;
    reg [7:0] z5141_assgn51410;
    reg [7:0] z5141_assgn51411;
    reg [7:0] z5141_assgn51412;
    reg [7:0] z2211_assgn2211;
    wire [7:0]  ny1_G256_newbasis1;
    wire [7:0]  z5145_assgn5145;
    reg [7:0] z5145_assgn51450;
    reg [7:0] z5145_assgn51451;
    reg [7:0] z5145_assgn51452;
    reg [7:0] z2214_assgn2214;
    wire [7:0]  tempybooloNegCond1_G256_newbasis1;
    wire [7:0]  y1_G256_newbasis1;
    wire [7:0]  z5151_assgn5151;
    reg [7:0] z5151_assgn51510;
    reg [7:0] z5151_assgn51511;
    reg [7:0] z5151_assgn51512;
    reg [7:0] z2217_assgn2217;
    wire [7:0]  x1_G256_newbasis1;
    wire [7:0]  tempy2_G256_newbasis1;
    wire [7:0]  z5157_assgn5157;
    reg [7:0] z5157_assgn51570;
    reg [7:0] z5157_assgn51571;
    reg [7:0] z5157_assgn51572;
    reg [7:0] z2221_assgn2221;
    wire [7:0]  cond2_G256_newbasis1;
    wire [7:0]  negCond2_G256_newbasis1;
    wire [7:0]  z5163_assgn5163;
    reg [7:0] z5163_assgn51630;
    reg [7:0] z5163_assgn51631;
    reg [7:0] z5163_assgn51632;
    reg [7:0] z2225_assgn2225;
    wire [7:0]  yxorb2_G256_newbasis1;
    wire [7:0]  ny2_G256_newbasis1;
    wire [7:0]  tempybooloNegCond2_G256_newbasis1;
    wire [7:0]  y2_G256_newbasis1;
    wire [7:0]  z5173_assgn5173;
    reg [7:0] z5173_assgn51730;
    reg [7:0] z5173_assgn51731;
    reg [7:0] z5173_assgn51732;
    reg [7:0] z2233_assgn2233;
    wire [7:0]  x2_G256_newbasis1;
    wire [7:0]  tempy3_G256_newbasis1;
    wire [7:0]  z5179_assgn5179;
    reg [7:0] z5179_assgn51790;
    reg [7:0] z5179_assgn51791;
    reg [7:0] z5179_assgn51792;
    reg [7:0] z2237_assgn2237;
    wire [7:0]  cond3_G256_newbasis1;
    wire [7:0]  negCond3_G256_newbasis1;
    wire [7:0]  z5185_assgn5185;
    reg [7:0] z5185_assgn51850;
    reg [7:0] z5185_assgn51851;
    reg [7:0] z5185_assgn51852;
    reg [7:0] z2241_assgn2241;
    wire [7:0]  yxorb3_G256_newbasis1;
    wire [7:0]  ny3_G256_newbasis1;
    wire [7:0]  tempybooloNegCond3_G256_newbasis1;
    wire [7:0]  y3_G256_newbasis1;
    wire [7:0]  z5195_assgn5195;
    reg [7:0] z5195_assgn51950;
    reg [7:0] z5195_assgn51951;
    reg [7:0] z5195_assgn51952;
    reg [7:0] z2249_assgn2249;
    wire [7:0]  x3_G256_newbasis1;
    wire [7:0]  tempy4_G256_newbasis1;
    wire [7:0]  z5201_assgn5201;
    reg [7:0] z5201_assgn52010;
    reg [7:0] z5201_assgn52011;
    reg [7:0] z5201_assgn52012;
    reg [7:0] z2253_assgn2253;
    wire [7:0]  cond4_G256_newbasis1;
    wire [7:0]  negCond4_G256_newbasis1;
    wire [7:0]  z5207_assgn5207;
    reg [7:0] z5207_assgn52070;
    reg [7:0] z5207_assgn52071;
    reg [7:0] z5207_assgn52072;
    reg [7:0] z2257_assgn2257;
    wire [7:0]  yxorb4_G256_newbasis1;
    wire [7:0]  ny4_G256_newbasis1;
    wire [7:0]  tempybooloNegCond4_G256_newbasis1;
    wire [7:0]  y4_G256_newbasis1;
    wire [7:0]  z5217_assgn5217;
    reg [7:0] z5217_assgn52170;
    reg [7:0] z5217_assgn52171;
    reg [7:0] z5217_assgn52172;
    reg [7:0] z2265_assgn2265;
    wire [7:0]  x4_G256_newbasis1;
    wire [7:0]  tempy5_G256_newbasis1;
    wire [7:0]  z5223_assgn5223;
    reg [7:0] z5223_assgn52230;
    reg [7:0] z5223_assgn52231;
    reg [7:0] z5223_assgn52232;
    reg [7:0] z2269_assgn2269;
    wire [7:0]  cond5_G256_newbasis1;
    wire [7:0]  negCond5_G256_newbasis1;
    wire [7:0]  z5229_assgn5229;
    reg [7:0] z5229_assgn52290;
    reg [7:0] z5229_assgn52291;
    reg [7:0] z5229_assgn52292;
    reg [7:0] z2273_assgn2273;
    wire [7:0]  yxorb5_G256_newbasis1;
    wire [7:0]  ny5_G256_newbasis1;
    wire [7:0]  tempybooloNegCond5_G256_newbasis1;
    wire [7:0]  y5_G256_newbasis1;
    wire [7:0]  z5239_assgn5239;
    reg [7:0] z5239_assgn52390;
    reg [7:0] z5239_assgn52391;
    reg [7:0] z5239_assgn52392;
    reg [7:0] z2281_assgn2281;
    wire [7:0]  x5_G256_newbasis1;
    wire [7:0]  tempy6_G256_newbasis1;
    wire [7:0]  z5245_assgn5245;
    reg [7:0] z5245_assgn52450;
    reg [7:0] z5245_assgn52451;
    reg [7:0] z5245_assgn52452;
    reg [7:0] z2285_assgn2285;
    wire [7:0]  cond6_G256_newbasis1;
    wire [7:0]  negCond6_G256_newbasis1;
    wire [7:0]  z5251_assgn5251;
    reg [7:0] z5251_assgn52510;
    reg [7:0] z5251_assgn52511;
    reg [7:0] z5251_assgn52512;
    reg [7:0] z2289_assgn2289;
    wire [7:0]  yxorb6_G256_newbasis1;
    wire [7:0]  ny6_G256_newbasis1;
    wire [7:0]  tempybooloNegCond6_G256_newbasis1;
    wire [7:0]  y6_G256_newbasis1;
    wire [7:0]  z5261_assgn5261;
    reg [7:0] z5261_assgn52610;
    reg [7:0] z5261_assgn52611;
    reg [7:0] z5261_assgn52612;
    reg [7:0] z2297_assgn2297;
    wire [7:0]  x6_G256_newbasis1;
    wire [7:0]  tempy7_G256_newbasis1;
    wire [7:0]  z5267_assgn5267;
    reg [7:0] z5267_assgn52670;
    reg [7:0] z5267_assgn52671;
    reg [7:0] z5267_assgn52672;
    reg [7:0] z2301_assgn2301;
    wire [7:0]  cond7_G256_newbasis1;
    wire [7:0]  negCond7_G256_newbasis1;
    wire [7:0]  z5273_assgn5273;
    reg [7:0] z5273_assgn52730;
    reg [7:0] z5273_assgn52731;
    reg [7:0] z5273_assgn52732;
    reg [7:0] z2305_assgn2305;
    wire [7:0]  yxorb7_G256_newbasis1;
    wire [7:0]  ny7_G256_newbasis1;
    wire [7:0]  tempybooloNegCond7_G256_newbasis1;
    wire [7:0]  y7_G256_newbasis1;
    wire [7:0]  z5283_assgn5283;
    reg [7:0] z5283_assgn52830;
    reg [7:0] z5283_assgn52831;
    reg [7:0] z5283_assgn52832;
    reg [7:0] z2313_assgn2313;
    wire [7:0]  x7_G256_newbasis1;
    wire [7:0]  tempy8_G256_newbasis1;
    wire [7:0]  z5289_assgn5289;
    reg [7:0] z5289_assgn52890;
    reg [7:0] z5289_assgn52891;
    reg [7:0] z5289_assgn52892;
    reg [7:0] z2317_assgn2317;
    wire [7:0]  cond8_G256_newbasis1;
    wire [7:0]  negCond8_G256_newbasis1;
    wire [7:0]  z5295_assgn5295;
    reg [7:0] z5295_assgn52950;
    reg [7:0] z5295_assgn52951;
    reg [7:0] z5295_assgn52952;
    reg [7:0] z2321_assgn2321;
    wire [7:0]  yxorb8_G256_newbasis1;
    wire [7:0]  ny8_G256_newbasis1;
    wire [7:0]  tempybooloNegCond8_G256_newbasis1;
    wire [7:0]  y8_G256_newbasis1;
    wire [7:0]  z5305_assgn5305;
    reg [7:0] z5305_assgn53050;
    reg [7:0] z5305_assgn53051;
    reg [7:0] z5305_assgn53052;
    reg [7:0] z2329_assgn2329;
    wire [7:0]  x8_G256_newbasis1;
    wire [7:0]  t6;
    wire [7:0]  z_y_G256_newbasis1;
    wire [7:0]  z_tempy1_G256_newbasis1;
    wire [7:0]  z5315_assgn5315;
    reg [7:0] z5315_assgn53150;
    reg [7:0] z5315_assgn53151;
    reg [7:0] z5315_assgn53152;
    reg [7:0] z2337_assgn2337;
    wire [7:0]  z_cond1_G256_newbasis1;
    wire [7:0]  z_negCond1_G256_newbasis1;
    wire [7:0]  z_yxorb1_G256_newbasis1;
    wire [7:0]  z5323_assgn5323;
    reg [7:0] z5323_assgn53230;
    reg [7:0] z5323_assgn53231;
    reg [7:0] z5323_assgn53232;
    reg [7:0] z2343_assgn2343;
    wire [7:0]  z_ny1_G256_newbasis1;
    wire [7:0]  z5327_assgn5327;
    reg [7:0] z5327_assgn53270;
    reg [7:0] z5327_assgn53271;
    reg [7:0] z5327_assgn53272;
    reg [7:0] z2346_assgn2346;
    wire [7:0]  z_tempybooloNegCond1_G256_newbasis1;
    wire [7:0]  z_y1_G256_newbasis1;
    wire [7:0]  z5333_assgn5333;
    reg [7:0] z5333_assgn53330;
    reg [7:0] z5333_assgn53331;
    reg [7:0] z5333_assgn53332;
    reg [7:0] z2349_assgn2349;
    wire [7:0]  z_x1_G256_newbasis1;
    wire [7:0]  z_tempy2_G256_newbasis1;
    wire [7:0]  z5339_assgn5339;
    reg [7:0] z5339_assgn53390;
    reg [7:0] z5339_assgn53391;
    reg [7:0] z5339_assgn53392;
    reg [7:0] z2353_assgn2353;
    wire [7:0]  z_cond2_G256_newbasis1;
    wire [7:0]  z_negCond2_G256_newbasis1;
    wire [7:0]  z5345_assgn5345;
    reg [7:0] z5345_assgn53450;
    reg [7:0] z5345_assgn53451;
    reg [7:0] z5345_assgn53452;
    reg [7:0] z2357_assgn2357;
    wire [7:0]  z_yxorb2_G256_newbasis1;
    wire [7:0]  z_ny2_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond2_G256_newbasis1;
    wire [7:0]  z_y2_G256_newbasis1;
    wire [7:0]  z5355_assgn5355;
    reg [7:0] z5355_assgn53550;
    reg [7:0] z5355_assgn53551;
    reg [7:0] z5355_assgn53552;
    reg [7:0] z2365_assgn2365;
    wire [7:0]  z_x2_G256_newbasis1;
    wire [7:0]  z_tempy3_G256_newbasis1;
    wire [7:0]  z5361_assgn5361;
    reg [7:0] z5361_assgn53610;
    reg [7:0] z5361_assgn53611;
    reg [7:0] z5361_assgn53612;
    reg [7:0] z2369_assgn2369;
    wire [7:0]  z_cond3_G256_newbasis1;
    wire [7:0]  z_negCond3_G256_newbasis1;
    wire [7:0]  z5367_assgn5367;
    reg [7:0] z5367_assgn53670;
    reg [7:0] z5367_assgn53671;
    reg [7:0] z5367_assgn53672;
    reg [7:0] z2373_assgn2373;
    wire [7:0]  z_yxorb3_G256_newbasis1;
    wire [7:0]  z_ny3_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond3_G256_newbasis1;
    wire [7:0]  z_y3_G256_newbasis1;
    wire [7:0]  z5377_assgn5377;
    reg [7:0] z5377_assgn53770;
    reg [7:0] z5377_assgn53771;
    reg [7:0] z5377_assgn53772;
    reg [7:0] z2381_assgn2381;
    wire [7:0]  z_x3_G256_newbasis1;
    wire [7:0]  z_tempy4_G256_newbasis1;
    wire [7:0]  z5383_assgn5383;
    reg [7:0] z5383_assgn53830;
    reg [7:0] z5383_assgn53831;
    reg [7:0] z5383_assgn53832;
    reg [7:0] z2385_assgn2385;
    wire [7:0]  z_cond4_G256_newbasis1;
    wire [7:0]  z_negCond4_G256_newbasis1;
    wire [7:0]  z5389_assgn5389;
    reg [7:0] z5389_assgn53890;
    reg [7:0] z5389_assgn53891;
    reg [7:0] z5389_assgn53892;
    reg [7:0] z2389_assgn2389;
    wire [7:0]  z_yxorb4_G256_newbasis1;
    wire [7:0]  z_ny4_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond4_G256_newbasis1;
    wire [7:0]  z_y4_G256_newbasis1;
    wire [7:0]  z5399_assgn5399;
    reg [7:0] z5399_assgn53990;
    reg [7:0] z5399_assgn53991;
    reg [7:0] z5399_assgn53992;
    reg [7:0] z2397_assgn2397;
    wire [7:0]  z_x4_G256_newbasis1;
    wire [7:0]  z_tempy5_G256_newbasis1;
    wire [7:0]  z5405_assgn5405;
    reg [7:0] z5405_assgn54050;
    reg [7:0] z5405_assgn54051;
    reg [7:0] z5405_assgn54052;
    reg [7:0] z2401_assgn2401;
    wire [7:0]  z_cond5_G256_newbasis1;
    wire [7:0]  z_negCond5_G256_newbasis1;
    wire [7:0]  z5411_assgn5411;
    reg [7:0] z5411_assgn54110;
    reg [7:0] z5411_assgn54111;
    reg [7:0] z5411_assgn54112;
    reg [7:0] z2405_assgn2405;
    wire [7:0]  z_yxorb5_G256_newbasis1;
    wire [7:0]  z_ny5_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond5_G256_newbasis1;
    wire [7:0]  z_y5_G256_newbasis1;
    wire [7:0]  z5421_assgn5421;
    reg [7:0] z5421_assgn54210;
    reg [7:0] z5421_assgn54211;
    reg [7:0] z5421_assgn54212;
    reg [7:0] z2413_assgn2413;
    wire [7:0]  z_x5_G256_newbasis1;
    wire [7:0]  z_tempy6_G256_newbasis1;
    wire [7:0]  z5427_assgn5427;
    reg [7:0] z5427_assgn54270;
    reg [7:0] z5427_assgn54271;
    reg [7:0] z5427_assgn54272;
    reg [7:0] z2417_assgn2417;
    wire [7:0]  z_cond6_G256_newbasis1;
    wire [7:0]  z_negCond6_G256_newbasis1;
    wire [7:0]  z5433_assgn5433;
    reg [7:0] z5433_assgn54330;
    reg [7:0] z5433_assgn54331;
    reg [7:0] z5433_assgn54332;
    reg [7:0] z2421_assgn2421;
    wire [7:0]  z_yxorb6_G256_newbasis1;
    wire [7:0]  z_ny6_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond6_G256_newbasis1;
    wire [7:0]  z_y6_G256_newbasis1;
    wire [7:0]  z5443_assgn5443;
    reg [7:0] z5443_assgn54430;
    reg [7:0] z5443_assgn54431;
    reg [7:0] z5443_assgn54432;
    reg [7:0] z2429_assgn2429;
    wire [7:0]  z_x6_G256_newbasis1;
    wire [7:0]  z_tempy7_G256_newbasis1;
    wire [7:0]  z5449_assgn5449;
    reg [7:0] z5449_assgn54490;
    reg [7:0] z5449_assgn54491;
    reg [7:0] z5449_assgn54492;
    reg [7:0] z2433_assgn2433;
    wire [7:0]  z_cond7_G256_newbasis1;
    wire [7:0]  z_negCond7_G256_newbasis1;
    wire [7:0]  z5455_assgn5455;
    reg [7:0] z5455_assgn54550;
    reg [7:0] z5455_assgn54551;
    reg [7:0] z5455_assgn54552;
    reg [7:0] z2437_assgn2437;
    wire [7:0]  z_yxorb7_G256_newbasis1;
    wire [7:0]  z_ny7_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond7_G256_newbasis1;
    wire [7:0]  z_y7_G256_newbasis1;
    wire [7:0]  z5465_assgn5465;
    reg [7:0] z5465_assgn54650;
    reg [7:0] z5465_assgn54651;
    reg [7:0] z5465_assgn54652;
    reg [7:0] z2445_assgn2445;
    wire [7:0]  z_x7_G256_newbasis1;
    wire [7:0]  z_tempy8_G256_newbasis1;
    wire [7:0]  z5471_assgn5471;
    reg [7:0] z5471_assgn54710;
    reg [7:0] z5471_assgn54711;
    reg [7:0] z5471_assgn54712;
    reg [7:0] z2449_assgn2449;
    wire [7:0]  z_cond8_G256_newbasis1;
    wire [7:0]  z_negCond8_G256_newbasis1;
    wire [7:0]  z5477_assgn5477;
    reg [7:0] z5477_assgn54770;
    reg [7:0] z5477_assgn54771;
    reg [7:0] z5477_assgn54772;
    reg [7:0] z2453_assgn2453;
    wire [7:0]  z_yxorb8_G256_newbasis1;
    wire [7:0]  z_ny8_G256_newbasis1;
    wire [7:0]  z_tempybooloNegCond8_G256_newbasis1;
    wire [7:0]  z_y8_G256_newbasis1;
    wire [7:0]  z5487_assgn5487;
    reg [7:0] z5487_assgn54870;
    reg [7:0] z5487_assgn54871;
    reg [7:0] z5487_assgn54872;
    reg [7:0] z2461_assgn2461;
    wire [7:0]  z_x8_G256_newbasis1;
    wire [7:0]  t7;
    wire [7:0]  z5493_assgn5493;
    reg [7:0] z5493_assgn54930;
    reg [7:0] z5493_assgn54931;
    reg [7:0] z5493_assgn54932;
    reg [7:0] z2465_assgn2465;

    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign r6_inp = r6;
    assign r7_inp = r7;
    assign r8_inp = r8;
    assign r9_inp = r9;
    assign r10_inp = r10;
    assign r11_inp = r11;
    assign r12_inp = r12;
    assign r13_inp = r13;
    assign r14_inp = r14;
    assign r15_inp = r15;
    assign r16_inp = r16;
    assign r17_inp = r17;
    assign r18_inp = r18;
    assign r19_inp = r19;
    assign r20_inp = r20;
    assign r21_inp = r21;
    assign r22_inp = r22;
    assign r23_inp = r23;
    assign r24_inp = r24;
    assign r25_inp = r25;
    assign r26_inp = r26;
    assign r27_inp = r27;
    assign r28_inp = r28;
    assign r29_inp = r29;
    assign r30_inp = r30;
    assign r31_inp = r31;
    assign r32_inp = r32;
    assign r33_inp = r33;
    assign r34_inp = r34;
    assign r35_inp = r35;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempybooloNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempybooloNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempybooloNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempybooloNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempybooloNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempybooloNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempybooloNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempybooloNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempybooloNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempybooloNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempybooloNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempybooloNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempybooloNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempybooloNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempybooloNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempybooloNegCond8_G256_newbasis0);
    assign z2721_assgn2721 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempybooloNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempybooloNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempybooloNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempybooloNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempybooloNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempybooloNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempybooloNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempybooloNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempybooloNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempybooloNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempybooloNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempybooloNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempybooloNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempybooloNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempybooloNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempybooloNegCond8_G256_newbasis0);
    assign z2853_assgn2853 = (z_x7_G256_newbasis0 >> dec_1_inp);
    assign t3 = z_y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a1_0_G256_inv0 = (t3 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a1xorb1_G256_inv0 = (a1_G256_inv0 ^ b1_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul0_G256_inv0 = (r5_inp % dec_16_inp);
    assign r60_G16_mul0_G256_inv0 = (r6_inp % dec_16_inp);
    assign r70_G16_mul0_G256_inv0 = (r7_inp % dec_16_inp);
    assign r80_G16_mul0_G256_inv0 = (r8_inp % dec_16_inp);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ d1_G4_mul0_G16_mul0_G256_inv0);
    assign z0_domand0_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 & cxord_1_G4_mul0_G16_mul0_G256_inv0);
    assign i1_domand0_G4_mul0_G16_mul0_G256_inv0 = (p2_domand0_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul0_G16_mul0_G256_inv0);
    assign p3_domand0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 & cxord_0_G4_mul0_G16_mul0_G256_inv0);
    assign i2_domand0_G4_mul0_G16_mul0_G256_inv0 = (p3_domand0_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_domand0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 & cxord_0_G4_mul0_G16_mul0_G256_inv0);
    assign p4_domand0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 & cxord_1_G4_mul0_G16_mul0_G256_inv0);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (i1_domand0_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_domand0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (i2_domand0_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_domand0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign z0_domand1_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 & c1_G4_mul0_G16_mul0_G256_inv0);
    assign i1_domand1_G4_mul0_G16_mul0_G256_inv0 = (p2_domand1_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul0_G16_mul0_G256_inv0);
    assign p3_domand1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 & c0_G4_mul0_G16_mul0_G256_inv0);
    assign i2_domand1_G4_mul0_G16_mul0_G256_inv0 = (p3_domand1_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul0_G16_mul0_G256_inv0);
    assign p1_domand1_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 & c0_G4_mul0_G16_mul0_G256_inv0);
    assign p4_domand1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 & c1_G4_mul0_G16_mul0_G256_inv0);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (i1_domand1_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_domand1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (i2_domand1_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_domand1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign z0_domand2_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 & d1_G4_mul0_G16_mul0_G256_inv0);
    assign i1_domand2_G4_mul0_G16_mul0_G256_inv0 = (p2_domand2_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul0_G16_mul0_G256_inv0);
    assign p3_domand2_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 & d0_G4_mul0_G16_mul0_G256_inv0);
    assign i2_domand2_G4_mul0_G16_mul0_G256_inv0 = (p3_domand2_G4_mul0_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul0_G16_mul0_G256_inv0);
    assign p1_domand2_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 & d0_G4_mul0_G16_mul0_G256_inv0);
    assign p4_domand2_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 & d1_G4_mul0_G16_mul0_G256_inv0);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (i1_domand2_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_domand2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (i2_domand2_G4_mul0_G16_mul0_G256_inv0_reg ^ p4_domand2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_2_inp_reg);
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & dec_2_inp_reg);
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp_reg);
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp_reg);
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_1_inp_reg);
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & dec_1_inp_reg);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ d1_G4_mul1_G16_mul0_G256_inv0);
    assign z0_domand0_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 & cxord_1_G4_mul1_G16_mul0_G256_inv0);
    assign i1_domand0_G4_mul1_G16_mul0_G256_inv0 = (p2_domand0_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul1_G16_mul0_G256_inv0);
    assign p3_domand0_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 & cxord_0_G4_mul1_G16_mul0_G256_inv0);
    assign i2_domand0_G4_mul1_G16_mul0_G256_inv0 = (p3_domand0_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_domand0_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 & cxord_0_G4_mul1_G16_mul0_G256_inv0);
    assign p4_domand0_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 & cxord_1_G4_mul1_G16_mul0_G256_inv0);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (i1_domand0_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_domand0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (i2_domand0_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_domand0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign z0_domand1_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 & c1_G4_mul1_G16_mul0_G256_inv0);
    assign i1_domand1_G4_mul1_G16_mul0_G256_inv0 = (p2_domand1_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul1_G16_mul0_G256_inv0);
    assign p3_domand1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 & c0_G4_mul1_G16_mul0_G256_inv0);
    assign i2_domand1_G4_mul1_G16_mul0_G256_inv0 = (p3_domand1_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_domand1_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 & c0_G4_mul1_G16_mul0_G256_inv0);
    assign p4_domand1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 & c1_G4_mul1_G16_mul0_G256_inv0);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (i1_domand1_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_domand1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (i2_domand1_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_domand1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign z0_domand2_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 & d1_G4_mul1_G16_mul0_G256_inv0);
    assign i1_domand2_G4_mul1_G16_mul0_G256_inv0 = (p2_domand2_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul1_G16_mul0_G256_inv0);
    assign p3_domand2_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 & d0_G4_mul1_G16_mul0_G256_inv0);
    assign i2_domand2_G4_mul1_G16_mul0_G256_inv0 = (p3_domand2_G4_mul1_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul1_G16_mul0_G256_inv0);
    assign p1_domand2_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 & d0_G4_mul1_G16_mul0_G256_inv0);
    assign p4_domand2_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 & d1_G4_mul1_G16_mul0_G256_inv0);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (i1_domand2_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_domand2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (i2_domand2_G4_mul1_G16_mul0_G256_inv0_reg ^ p4_domand2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r60_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r70_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r80_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ d1_G4_mul2_G16_mul0_G256_inv0);
    assign z0_domand0_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 & cxord_1_G4_mul2_G16_mul0_G256_inv0);
    assign i1_domand0_G4_mul2_G16_mul0_G256_inv0 = (p2_domand0_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul2_G16_mul0_G256_inv0);
    assign p3_domand0_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 & cxord_0_G4_mul2_G16_mul0_G256_inv0);
    assign i2_domand0_G4_mul2_G16_mul0_G256_inv0 = (p3_domand0_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_domand0_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 & cxord_0_G4_mul2_G16_mul0_G256_inv0);
    assign p4_domand0_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 & cxord_1_G4_mul2_G16_mul0_G256_inv0);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (i1_domand0_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_domand0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (i2_domand0_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_domand0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign z0_domand1_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 & c1_G4_mul2_G16_mul0_G256_inv0);
    assign i1_domand1_G4_mul2_G16_mul0_G256_inv0 = (p2_domand1_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul2_G16_mul0_G256_inv0);
    assign p3_domand1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 & c0_G4_mul2_G16_mul0_G256_inv0);
    assign i2_domand1_G4_mul2_G16_mul0_G256_inv0 = (p3_domand1_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand1_G4_mul2_G16_mul0_G256_inv0);
    assign p1_domand1_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 & c0_G4_mul2_G16_mul0_G256_inv0);
    assign p4_domand1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 & c1_G4_mul2_G16_mul0_G256_inv0);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (i1_domand1_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_domand1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (i2_domand1_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_domand1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign z0_domand2_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 & d1_G4_mul2_G16_mul0_G256_inv0);
    assign i1_domand2_G4_mul2_G16_mul0_G256_inv0 = (p2_domand2_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul2_G16_mul0_G256_inv0);
    assign p3_domand2_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 & d0_G4_mul2_G16_mul0_G256_inv0);
    assign i2_domand2_G4_mul2_G16_mul0_G256_inv0 = (p3_domand2_G4_mul2_G16_mul0_G256_inv0 ^ z0_domand2_G4_mul2_G16_mul0_G256_inv0);
    assign p1_domand2_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 & d0_G4_mul2_G16_mul0_G256_inv0);
    assign p4_domand2_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 & d1_G4_mul2_G16_mul0_G256_inv0);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (i1_domand2_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_domand2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (i2_domand2_G4_mul2_G16_mul0_G256_inv0_reg ^ p4_domand2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp_reg);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << dec_2_inp_reg);
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << dec_2_inp_reg);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign c0xord0_G256_inv0 = (c0_G256_inv0_reg ^ d0_G256_inv0);
    assign c1xord1_G256_inv0 = (c1_G256_inv0_reg ^ d1_G256_inv0);
    assign r00_G16_inv0_G256_inv0 = (r9_inp % dec_16_inp);
    assign r10_G16_inv0_G256_inv0 = (r10_inp % dec_16_inp);
    assign r20_G16_inv0_G256_inv0 = (r11_inp % dec_16_inp);
    assign r30_G16_inv0_G256_inv0 = (r12_inp % dec_16_inp);
    assign r40_G16_inv0_G256_inv0 = (r13_inp % dec_16_inp);
    assign r50_G16_inv0_G256_inv0 = (r14_inp % dec_16_inp);
    assign r60_G16_inv0_G256_inv0 = (r15_inp % dec_16_inp);
    assign r70_G16_inv0_G256_inv0 = (r16_inp % dec_16_inp);
    assign r80_G16_inv0_G256_inv0 = (r17_inp % dec_16_inp);
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_12_inp_reg);
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & dec_12_inp_reg);
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> dec_2_inp_reg);
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> dec_2_inp_reg);
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_3_inp_reg);
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & dec_3_inp_reg);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a1xorb1_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 ^ b1_G16_inv0_G256_inv0);
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp_reg);
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp_reg);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp_reg);
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp_reg);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ d1_G4_mul3_G16_inv0_G256_inv0);
    assign z0_domand0_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 & cxord_1_G4_mul3_G16_inv0_G256_inv0);
    assign i1_domand0_G4_mul3_G16_inv0_G256_inv0 = (p2_domand0_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_domand0_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 & cxord_0_G4_mul3_G16_inv0_G256_inv0);
    assign i2_domand0_G4_mul3_G16_inv0_G256_inv0 = (p3_domand0_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_domand0_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 & cxord_0_G4_mul3_G16_inv0_G256_inv0);
    assign p4_domand0_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 & cxord_1_G4_mul3_G16_inv0_G256_inv0);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (i1_domand0_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_domand0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (i2_domand0_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_domand0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z0_domand1_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 & c1_G4_mul3_G16_inv0_G256_inv0);
    assign i1_domand1_G4_mul3_G16_inv0_G256_inv0 = (p2_domand1_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_domand1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 & c0_G4_mul3_G16_inv0_G256_inv0);
    assign i2_domand1_G4_mul3_G16_inv0_G256_inv0 = (p3_domand1_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_domand1_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 & c0_G4_mul3_G16_inv0_G256_inv0);
    assign p4_domand1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 & c1_G4_mul3_G16_inv0_G256_inv0);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (i1_domand1_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_domand1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (i2_domand1_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_domand1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z0_domand2_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 & d1_G4_mul3_G16_inv0_G256_inv0);
    assign i1_domand2_G4_mul3_G16_inv0_G256_inv0 = (p2_domand2_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_domand2_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 & d0_G4_mul3_G16_inv0_G256_inv0);
    assign i2_domand2_G4_mul3_G16_inv0_G256_inv0 = (p3_domand2_G4_mul3_G16_inv0_G256_inv0 ^ z0_domand2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_domand2_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 & d0_G4_mul3_G16_inv0_G256_inv0);
    assign p4_domand2_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 & d1_G4_mul3_G16_inv0_G256_inv0);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (i1_domand2_G4_mul3_G16_inv0_G256_inv0_reg ^ p1_domand2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (i2_domand2_G4_mul3_G16_inv0_G256_inv0_reg ^ p4_domand2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z3569_assgn3569 = dec_1_inp;
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << z1101_assgn1101);
    assign z3573_assgn3573 = dec_1_inp;
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << z1103_assgn1103);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign c0xord0_G16_inv0_G256_inv0 = (c0_G16_inv0_G256_inv0_reg ^ d0_G16_inv0_G256_inv0);
    assign c1xord1_G16_inv0_G256_inv0 = (c1_G16_inv0_G256_inv0_reg ^ d1_G16_inv0_G256_inv0);
    assign z3585_assgn3585 = dec_2_inp;
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1113_assgn1113);
    assign z3589_assgn3589 = dec_2_inp;
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1115_assgn1115);
    assign z3593_assgn3593 = dec_1_inp;
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> z1117_assgn1117);
    assign z3597_assgn3597 = dec_1_inp;
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> z1119_assgn1119);
    assign z3601_assgn3601 = dec_1_inp;
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1121_assgn1121);
    assign z3605_assgn3605 = dec_1_inp;
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1123_assgn1123);
    assign z3609_assgn3609 = dec_1_inp;
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << z1125_assgn1125);
    assign z3613_assgn3613 = dec_1_inp;
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << z1127_assgn1127);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign z3627_assgn3627 = dec_2_inp;
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1139_assgn1139);
    assign z3631_assgn3631 = dec_2_inp;
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1141_assgn1141);
    assign z3635_assgn3635 = dec_1_inp;
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> z1143_assgn1143);
    assign z3639_assgn3639 = dec_1_inp;
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> z1145_assgn1145);
    assign z3643_assgn3643 = dec_1_inp;
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1147_assgn1147);
    assign z3647_assgn3647 = dec_1_inp;
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1149_assgn1149);
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ d1_G4_mul4_G16_inv0_G256_inv0);
    assign z0_domand0_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & cxord_1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3675_assgn3675 = z0_domand0_G4_mul4_G16_inv0_G256_inv0;
    assign i1_domand0_G4_mul4_G16_inv0_G256_inv0 = (p2_domand0_G4_mul4_G16_inv0_G256_inv0 ^ z1175_assgn1175);
    assign p3_domand0_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & cxord_0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3681_assgn3681 = z0_domand0_G4_mul4_G16_inv0_G256_inv0;
    assign i2_domand0_G4_mul4_G16_inv0_G256_inv0 = (p3_domand0_G4_mul4_G16_inv0_G256_inv0 ^ z1179_assgn1179);
    assign p1_domand0_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & cxord_0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p4_domand0_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & cxord_1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (i1_domand0_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_domand0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (i2_domand0_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_domand0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z0_domand1_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & c1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3697_assgn3697 = z0_domand1_G4_mul4_G16_inv0_G256_inv0;
    assign i1_domand1_G4_mul4_G16_inv0_G256_inv0 = (p2_domand1_G4_mul4_G16_inv0_G256_inv0 ^ z1193_assgn1193);
    assign p3_domand1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & c0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3703_assgn3703 = z0_domand1_G4_mul4_G16_inv0_G256_inv0;
    assign i2_domand1_G4_mul4_G16_inv0_G256_inv0 = (p3_domand1_G4_mul4_G16_inv0_G256_inv0 ^ z1197_assgn1197);
    assign p1_domand1_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & c0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p4_domand1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & c1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (i1_domand1_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_domand1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (i2_domand1_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_domand1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z0_domand2_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & d1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3723_assgn3723 = z0_domand2_G4_mul4_G16_inv0_G256_inv0;
    assign i1_domand2_G4_mul4_G16_inv0_G256_inv0 = (p2_domand2_G4_mul4_G16_inv0_G256_inv0 ^ z1215_assgn1215);
    assign p3_domand2_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & d0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z3729_assgn3729 = z0_domand2_G4_mul4_G16_inv0_G256_inv0;
    assign i2_domand2_G4_mul4_G16_inv0_G256_inv0 = (p3_domand2_G4_mul4_G16_inv0_G256_inv0 ^ z1219_assgn1219);
    assign p1_domand2_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & d0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p4_domand2_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & d1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (i1_domand2_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_domand2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (i2_domand2_G4_mul4_G16_inv0_G256_inv0_reg ^ p4_domand2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z3745_assgn3745 = dec_1_inp;
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << z1233_assgn1233);
    assign z3749_assgn3749 = dec_1_inp;
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << z1235_assgn1235);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r60_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r70_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r80_G16_inv0_G256_inv0 % dec_4_inp);
    assign z3763_assgn3763 = dec_2_inp;
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1247_assgn1247);
    assign z3767_assgn3767 = dec_2_inp;
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1249_assgn1249);
    assign z3771_assgn3771 = dec_1_inp;
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> z1251_assgn1251);
    assign z3775_assgn3775 = dec_1_inp;
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> z1253_assgn1253);
    assign z3779_assgn3779 = dec_1_inp;
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1255_assgn1255);
    assign z3783_assgn3783 = dec_1_inp;
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1257_assgn1257);
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_2_inp_reg);
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp_reg);
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_1_inp_reg);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ d1_G4_mul5_G16_inv0_G256_inv0);
    assign z0_domand0_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand0_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & cxord_1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3811_assgn3811 = z0_domand0_G4_mul5_G16_inv0_G256_inv0;
    assign i1_domand0_G4_mul5_G16_inv0_G256_inv0 = (p2_domand0_G4_mul5_G16_inv0_G256_inv0 ^ z1283_assgn1283);
    assign p3_domand0_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & cxord_0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3817_assgn3817 = z0_domand0_G4_mul5_G16_inv0_G256_inv0;
    assign i2_domand0_G4_mul5_G16_inv0_G256_inv0 = (p3_domand0_G4_mul5_G16_inv0_G256_inv0 ^ z1287_assgn1287);
    assign p1_domand0_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & cxord_0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p4_domand0_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & cxord_1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (i1_domand0_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_domand0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (i2_domand0_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_domand0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z0_domand1_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand1_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & c1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3833_assgn3833 = z0_domand1_G4_mul5_G16_inv0_G256_inv0;
    assign i1_domand1_G4_mul5_G16_inv0_G256_inv0 = (p2_domand1_G4_mul5_G16_inv0_G256_inv0 ^ z1301_assgn1301);
    assign p3_domand1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & c0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3839_assgn3839 = z0_domand1_G4_mul5_G16_inv0_G256_inv0;
    assign i2_domand1_G4_mul5_G16_inv0_G256_inv0 = (p3_domand1_G4_mul5_G16_inv0_G256_inv0 ^ z1305_assgn1305);
    assign p1_domand1_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & c0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p4_domand1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & c1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (i1_domand1_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_domand1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (i2_domand1_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_domand1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z0_domand2_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign p2_domand2_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & d1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3859_assgn3859 = z0_domand2_G4_mul5_G16_inv0_G256_inv0;
    assign i1_domand2_G4_mul5_G16_inv0_G256_inv0 = (p2_domand2_G4_mul5_G16_inv0_G256_inv0 ^ z1323_assgn1323);
    assign p3_domand2_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & d0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z3865_assgn3865 = z0_domand2_G4_mul5_G16_inv0_G256_inv0;
    assign i2_domand2_G4_mul5_G16_inv0_G256_inv0 = (p3_domand2_G4_mul5_G16_inv0_G256_inv0 ^ z1327_assgn1327);
    assign p1_domand2_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & d0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p4_domand2_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & d1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (i1_domand2_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_domand2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (i2_domand2_G4_mul5_G16_inv0_G256_inv0_reg ^ p4_domand2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z3881_assgn3881 = dec_1_inp;
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << z1341_assgn1341);
    assign z3885_assgn3885 = dec_1_inp;
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << z1343_assgn1343);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign z3893_assgn3893 = dec_2_inp;
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << z1349_assgn1349);
    assign z3897_assgn3897 = dec_2_inp;
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << z1351_assgn1351);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign r00_G16_mul1_G256_inv0 = (r18_inp % dec_16_inp);
    assign r10_G16_mul1_G256_inv0 = (r19_inp % dec_16_inp);
    assign r20_G16_mul1_G256_inv0 = (r20_inp % dec_16_inp);
    assign r30_G16_mul1_G256_inv0 = (r21_inp % dec_16_inp);
    assign r40_G16_mul1_G256_inv0 = (r22_inp % dec_16_inp);
    assign r50_G16_mul1_G256_inv0 = (r23_inp % dec_16_inp);
    assign r60_G16_mul1_G256_inv0 = (r24_inp % dec_16_inp);
    assign r70_G16_mul1_G256_inv0 = (r25_inp % dec_16_inp);
    assign r80_G16_mul1_G256_inv0 = (r26_inp % dec_16_inp);
    assign z3923_assgn3923 = dec_12_inp;
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1375_assgn1375);
    assign z3927_assgn3927 = dec_12_inp;
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1377_assgn1377);
    assign z3931_assgn3931 = dec_2_inp;
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> z1379_assgn1379);
    assign z3935_assgn3935 = dec_2_inp;
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> z1381_assgn1381);
    assign z3939_assgn3939 = dec_3_inp;
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1383_assgn1383);
    assign z3943_assgn3943 = dec_3_inp;
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1385_assgn1385);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign z3973_assgn3973 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1413_assgn1413);
    assign z3977_assgn3977 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1415_assgn1415);
    assign z3981_assgn3981 = dec_1_inp;
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> z1417_assgn1417);
    assign z3985_assgn3985 = dec_1_inp;
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> z1419_assgn1419);
    assign z3989_assgn3989 = dec_1_inp;
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1421_assgn1421);
    assign z3993_assgn3993 = dec_1_inp;
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1423_assgn1423);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ d1_G4_mul0_G16_mul1_G256_inv0);
    assign z0_domand0_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4019_assgn4019 = cxord_1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_domand0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1447_assgn1447);
    assign z4023_assgn4023 = z0_domand0_G4_mul0_G16_mul1_G256_inv0;
    assign i1_domand0_G4_mul0_G16_mul1_G256_inv0 = (p2_domand0_G4_mul0_G16_mul1_G256_inv0 ^ z1449_assgn1449);
    assign z4027_assgn4027 = cxord_0_G4_mul0_G16_mul1_G256_inv0;
    assign p3_domand0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1451_assgn1451);
    assign z4031_assgn4031 = z0_domand0_G4_mul0_G16_mul1_G256_inv0;
    assign i2_domand0_G4_mul0_G16_mul1_G256_inv0 = (p3_domand0_G4_mul0_G16_mul1_G256_inv0 ^ z1453_assgn1453);
    assign z4035_assgn4035 = cxord_0_G4_mul0_G16_mul1_G256_inv0;
    assign p1_domand0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1455_assgn1455);
    assign z4039_assgn4039 = cxord_1_G4_mul0_G16_mul1_G256_inv0;
    assign p4_domand0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1457_assgn1457);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (i1_domand0_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_domand0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (i2_domand0_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_domand0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z0_domand1_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4049_assgn4049 = c1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_domand1_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1465_assgn1465);
    assign z4053_assgn4053 = z0_domand1_G4_mul0_G16_mul1_G256_inv0;
    assign i1_domand1_G4_mul0_G16_mul1_G256_inv0 = (p2_domand1_G4_mul0_G16_mul1_G256_inv0 ^ z1467_assgn1467);
    assign z4057_assgn4057 = c0_G4_mul0_G16_mul1_G256_inv0;
    assign p3_domand1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1469_assgn1469);
    assign z4061_assgn4061 = z0_domand1_G4_mul0_G16_mul1_G256_inv0;
    assign i2_domand1_G4_mul0_G16_mul1_G256_inv0 = (p3_domand1_G4_mul0_G16_mul1_G256_inv0 ^ z1471_assgn1471);
    assign z4065_assgn4065 = c0_G4_mul0_G16_mul1_G256_inv0;
    assign p1_domand1_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1473_assgn1473);
    assign z4069_assgn4069 = c1_G4_mul0_G16_mul1_G256_inv0;
    assign p4_domand1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1475_assgn1475);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (i1_domand1_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_domand1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (i2_domand1_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_domand1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z0_domand2_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4083_assgn4083 = d1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_domand2_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1487_assgn1487);
    assign z4087_assgn4087 = z0_domand2_G4_mul0_G16_mul1_G256_inv0;
    assign i1_domand2_G4_mul0_G16_mul1_G256_inv0 = (p2_domand2_G4_mul0_G16_mul1_G256_inv0 ^ z1489_assgn1489);
    assign z4091_assgn4091 = d0_G4_mul0_G16_mul1_G256_inv0;
    assign p3_domand2_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1491_assgn1491);
    assign z4095_assgn4095 = z0_domand2_G4_mul0_G16_mul1_G256_inv0;
    assign i2_domand2_G4_mul0_G16_mul1_G256_inv0 = (p3_domand2_G4_mul0_G16_mul1_G256_inv0 ^ z1493_assgn1493);
    assign z4099_assgn4099 = d0_G4_mul0_G16_mul1_G256_inv0;
    assign p1_domand2_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1495_assgn1495);
    assign z4103_assgn4103 = d1_G4_mul0_G16_mul1_G256_inv0;
    assign p4_domand2_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1497_assgn1497);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (i1_domand2_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_domand2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (i2_domand2_G4_mul0_G16_mul1_G256_inv0_reg ^ p4_domand2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z4115_assgn4115 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << z1507_assgn1507);
    assign z4119_assgn4119 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << z1509_assgn1509);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign z4127_assgn4127 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1515_assgn1515);
    assign z4131_assgn4131 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1517_assgn1517);
    assign z4135_assgn4135 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1519_assgn1519);
    assign z4139_assgn4139 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1521_assgn1521);
    assign z4143_assgn4143 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1523_assgn1523);
    assign z4147_assgn4147 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1525_assgn1525);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z4159_assgn4159 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << z1535_assgn1535);
    assign z4163_assgn4163 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << z1537_assgn1537);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign z4177_assgn4177 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1549_assgn1549);
    assign z4181_assgn4181 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1551_assgn1551);
    assign z4185_assgn4185 = dec_1_inp;
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> z1553_assgn1553);
    assign z4189_assgn4189 = dec_1_inp;
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> z1555_assgn1555);
    assign z4193_assgn4193 = dec_1_inp;
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1557_assgn1557);
    assign z4197_assgn4197 = dec_1_inp;
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1559_assgn1559);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ d1_G4_mul1_G16_mul1_G256_inv0);
    assign z0_domand0_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4223_assgn4223 = cxord_1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_domand0_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1583_assgn1583);
    assign z4227_assgn4227 = z0_domand0_G4_mul1_G16_mul1_G256_inv0;
    assign i1_domand0_G4_mul1_G16_mul1_G256_inv0 = (p2_domand0_G4_mul1_G16_mul1_G256_inv0 ^ z1585_assgn1585);
    assign z4231_assgn4231 = cxord_0_G4_mul1_G16_mul1_G256_inv0;
    assign p3_domand0_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1587_assgn1587);
    assign z4235_assgn4235 = z0_domand0_G4_mul1_G16_mul1_G256_inv0;
    assign i2_domand0_G4_mul1_G16_mul1_G256_inv0 = (p3_domand0_G4_mul1_G16_mul1_G256_inv0 ^ z1589_assgn1589);
    assign z4239_assgn4239 = cxord_0_G4_mul1_G16_mul1_G256_inv0;
    assign p1_domand0_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1591_assgn1591);
    assign z4243_assgn4243 = cxord_1_G4_mul1_G16_mul1_G256_inv0;
    assign p4_domand0_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1593_assgn1593);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (i1_domand0_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_domand0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (i2_domand0_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_domand0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z0_domand1_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4253_assgn4253 = c1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_domand1_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1601_assgn1601);
    assign z4257_assgn4257 = z0_domand1_G4_mul1_G16_mul1_G256_inv0;
    assign i1_domand1_G4_mul1_G16_mul1_G256_inv0 = (p2_domand1_G4_mul1_G16_mul1_G256_inv0 ^ z1603_assgn1603);
    assign z4261_assgn4261 = c0_G4_mul1_G16_mul1_G256_inv0;
    assign p3_domand1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1605_assgn1605);
    assign z4265_assgn4265 = z0_domand1_G4_mul1_G16_mul1_G256_inv0;
    assign i2_domand1_G4_mul1_G16_mul1_G256_inv0 = (p3_domand1_G4_mul1_G16_mul1_G256_inv0 ^ z1607_assgn1607);
    assign z4269_assgn4269 = c0_G4_mul1_G16_mul1_G256_inv0;
    assign p1_domand1_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1609_assgn1609);
    assign z4273_assgn4273 = c1_G4_mul1_G16_mul1_G256_inv0;
    assign p4_domand1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1611_assgn1611);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (i1_domand1_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_domand1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (i2_domand1_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_domand1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z0_domand2_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4287_assgn4287 = d1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_domand2_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1623_assgn1623);
    assign z4291_assgn4291 = z0_domand2_G4_mul1_G16_mul1_G256_inv0;
    assign i1_domand2_G4_mul1_G16_mul1_G256_inv0 = (p2_domand2_G4_mul1_G16_mul1_G256_inv0 ^ z1625_assgn1625);
    assign z4295_assgn4295 = d0_G4_mul1_G16_mul1_G256_inv0;
    assign p3_domand2_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1627_assgn1627);
    assign z4299_assgn4299 = z0_domand2_G4_mul1_G16_mul1_G256_inv0;
    assign i2_domand2_G4_mul1_G16_mul1_G256_inv0 = (p3_domand2_G4_mul1_G16_mul1_G256_inv0 ^ z1629_assgn1629);
    assign z4303_assgn4303 = d0_G4_mul1_G16_mul1_G256_inv0;
    assign p1_domand2_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1631_assgn1631);
    assign z4307_assgn4307 = d1_G4_mul1_G16_mul1_G256_inv0;
    assign p4_domand2_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1633_assgn1633);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (i1_domand2_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_domand2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (i2_domand2_G4_mul1_G16_mul1_G256_inv0_reg ^ p4_domand2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z4319_assgn4319 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << z1643_assgn1643);
    assign z4323_assgn4323 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << z1645_assgn1645);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r60_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r70_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r80_G16_mul1_G256_inv0 % dec_4_inp);
    assign z4341_assgn4341 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1661_assgn1661);
    assign z4345_assgn4345 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1663_assgn1663);
    assign z4349_assgn4349 = dec_1_inp;
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> z1665_assgn1665);
    assign z4353_assgn4353 = dec_1_inp;
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> z1667_assgn1667);
    assign z4357_assgn4357 = dec_1_inp;
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1669_assgn1669);
    assign z4361_assgn4361 = dec_1_inp;
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1671_assgn1671);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ d1_G4_mul2_G16_mul1_G256_inv0);
    assign z0_domand0_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4387_assgn4387 = cxord_1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_domand0_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z1695_assgn1695);
    assign z4391_assgn4391 = z0_domand0_G4_mul2_G16_mul1_G256_inv0;
    assign i1_domand0_G4_mul2_G16_mul1_G256_inv0 = (p2_domand0_G4_mul2_G16_mul1_G256_inv0 ^ z1697_assgn1697);
    assign z4395_assgn4395 = cxord_0_G4_mul2_G16_mul1_G256_inv0;
    assign p3_domand0_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z1699_assgn1699);
    assign z4399_assgn4399 = z0_domand0_G4_mul2_G16_mul1_G256_inv0;
    assign i2_domand0_G4_mul2_G16_mul1_G256_inv0 = (p3_domand0_G4_mul2_G16_mul1_G256_inv0 ^ z1701_assgn1701);
    assign z4403_assgn4403 = cxord_0_G4_mul2_G16_mul1_G256_inv0;
    assign p1_domand0_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z1703_assgn1703);
    assign z4407_assgn4407 = cxord_1_G4_mul2_G16_mul1_G256_inv0;
    assign p4_domand0_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z1705_assgn1705);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (i1_domand0_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_domand0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (i2_domand0_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_domand0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z0_domand1_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4417_assgn4417 = c1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_domand1_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z1713_assgn1713);
    assign z4421_assgn4421 = z0_domand1_G4_mul2_G16_mul1_G256_inv0;
    assign i1_domand1_G4_mul2_G16_mul1_G256_inv0 = (p2_domand1_G4_mul2_G16_mul1_G256_inv0 ^ z1715_assgn1715);
    assign z4425_assgn4425 = c0_G4_mul2_G16_mul1_G256_inv0;
    assign p3_domand1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z1717_assgn1717);
    assign z4429_assgn4429 = z0_domand1_G4_mul2_G16_mul1_G256_inv0;
    assign i2_domand1_G4_mul2_G16_mul1_G256_inv0 = (p3_domand1_G4_mul2_G16_mul1_G256_inv0 ^ z1719_assgn1719);
    assign z4433_assgn4433 = c0_G4_mul2_G16_mul1_G256_inv0;
    assign p1_domand1_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z1721_assgn1721);
    assign z4437_assgn4437 = c1_G4_mul2_G16_mul1_G256_inv0;
    assign p4_domand1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z1723_assgn1723);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (i1_domand1_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_domand1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (i2_domand1_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_domand1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z0_domand2_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign z4451_assgn4451 = d1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_domand2_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z1735_assgn1735);
    assign z4455_assgn4455 = z0_domand2_G4_mul2_G16_mul1_G256_inv0;
    assign i1_domand2_G4_mul2_G16_mul1_G256_inv0 = (p2_domand2_G4_mul2_G16_mul1_G256_inv0 ^ z1737_assgn1737);
    assign z4459_assgn4459 = d0_G4_mul2_G16_mul1_G256_inv0;
    assign p3_domand2_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z1739_assgn1739);
    assign z4463_assgn4463 = z0_domand2_G4_mul2_G16_mul1_G256_inv0;
    assign i2_domand2_G4_mul2_G16_mul1_G256_inv0 = (p3_domand2_G4_mul2_G16_mul1_G256_inv0 ^ z1741_assgn1741);
    assign z4467_assgn4467 = d0_G4_mul2_G16_mul1_G256_inv0;
    assign p1_domand2_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z1743_assgn1743);
    assign z4471_assgn4471 = d1_G4_mul2_G16_mul1_G256_inv0;
    assign p4_domand2_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z1745_assgn1745);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (i1_domand2_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_domand2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (i2_domand2_G4_mul2_G16_mul1_G256_inv0_reg ^ p4_domand2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z4483_assgn4483 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << z1755_assgn1755);
    assign z4487_assgn4487 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << z1757_assgn1757);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign z4499_assgn4499 = dec_2_inp;
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << z1767_assgn1767);
    assign z4503_assgn4503 = dec_2_inp;
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << z1769_assgn1769);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign r00_G16_mul2_G256_inv0 = (r27_inp % dec_16_inp);
    assign r10_G16_mul2_G256_inv0 = (r28_inp % dec_16_inp);
    assign r20_G16_mul2_G256_inv0 = (r29_inp % dec_16_inp);
    assign r30_G16_mul2_G256_inv0 = (r30_inp % dec_16_inp);
    assign r40_G16_mul2_G256_inv0 = (r31_inp % dec_16_inp);
    assign r50_G16_mul2_G256_inv0 = (r32_inp % dec_16_inp);
    assign r60_G16_mul2_G256_inv0 = (r33_inp % dec_16_inp);
    assign r70_G16_mul2_G256_inv0 = (r34_inp % dec_16_inp);
    assign r80_G16_mul2_G256_inv0 = (r35_inp % dec_16_inp);
    assign z4529_assgn4529 = dec_12_inp;
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z1793_assgn1793);
    assign z4533_assgn4533 = dec_12_inp;
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & z1795_assgn1795);
    assign z4537_assgn4537 = dec_2_inp;
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> z1797_assgn1797);
    assign z4541_assgn4541 = dec_2_inp;
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> z1799_assgn1799);
    assign z4545_assgn4545 = dec_3_inp;
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z1801_assgn1801);
    assign z4549_assgn4549 = dec_3_inp;
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & z1803_assgn1803);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign z4579_assgn4579 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z1831_assgn1831);
    assign z4583_assgn4583 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z1833_assgn1833);
    assign z4587_assgn4587 = dec_1_inp;
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> z1835_assgn1835);
    assign z4591_assgn4591 = dec_1_inp;
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> z1837_assgn1837);
    assign z4595_assgn4595 = dec_1_inp;
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z1839_assgn1839);
    assign z4599_assgn4599 = dec_1_inp;
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z1841_assgn1841);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ d1_G4_mul0_G16_mul2_G256_inv0);
    assign z0_domand0_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4625_assgn4625 = cxord_1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_domand0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z1865_assgn1865);
    assign z4629_assgn4629 = z0_domand0_G4_mul0_G16_mul2_G256_inv0;
    assign i1_domand0_G4_mul0_G16_mul2_G256_inv0 = (p2_domand0_G4_mul0_G16_mul2_G256_inv0 ^ z1867_assgn1867);
    assign z4633_assgn4633 = cxord_0_G4_mul0_G16_mul2_G256_inv0;
    assign p3_domand0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z1869_assgn1869);
    assign z4637_assgn4637 = z0_domand0_G4_mul0_G16_mul2_G256_inv0;
    assign i2_domand0_G4_mul0_G16_mul2_G256_inv0 = (p3_domand0_G4_mul0_G16_mul2_G256_inv0 ^ z1871_assgn1871);
    assign z4641_assgn4641 = cxord_0_G4_mul0_G16_mul2_G256_inv0;
    assign p1_domand0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z1873_assgn1873);
    assign z4645_assgn4645 = cxord_1_G4_mul0_G16_mul2_G256_inv0;
    assign p4_domand0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z1875_assgn1875);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (i1_domand0_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_domand0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (i2_domand0_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_domand0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z0_domand1_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4655_assgn4655 = c1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_domand1_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z1883_assgn1883);
    assign z4659_assgn4659 = z0_domand1_G4_mul0_G16_mul2_G256_inv0;
    assign i1_domand1_G4_mul0_G16_mul2_G256_inv0 = (p2_domand1_G4_mul0_G16_mul2_G256_inv0 ^ z1885_assgn1885);
    assign z4663_assgn4663 = c0_G4_mul0_G16_mul2_G256_inv0;
    assign p3_domand1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z1887_assgn1887);
    assign z4667_assgn4667 = z0_domand1_G4_mul0_G16_mul2_G256_inv0;
    assign i2_domand1_G4_mul0_G16_mul2_G256_inv0 = (p3_domand1_G4_mul0_G16_mul2_G256_inv0 ^ z1889_assgn1889);
    assign z4671_assgn4671 = c0_G4_mul0_G16_mul2_G256_inv0;
    assign p1_domand1_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z1891_assgn1891);
    assign z4675_assgn4675 = c1_G4_mul0_G16_mul2_G256_inv0;
    assign p4_domand1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z1893_assgn1893);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (i1_domand1_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_domand1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (i2_domand1_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_domand1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z0_domand2_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4689_assgn4689 = d1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_domand2_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z1905_assgn1905);
    assign z4693_assgn4693 = z0_domand2_G4_mul0_G16_mul2_G256_inv0;
    assign i1_domand2_G4_mul0_G16_mul2_G256_inv0 = (p2_domand2_G4_mul0_G16_mul2_G256_inv0 ^ z1907_assgn1907);
    assign z4697_assgn4697 = d0_G4_mul0_G16_mul2_G256_inv0;
    assign p3_domand2_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z1909_assgn1909);
    assign z4701_assgn4701 = z0_domand2_G4_mul0_G16_mul2_G256_inv0;
    assign i2_domand2_G4_mul0_G16_mul2_G256_inv0 = (p3_domand2_G4_mul0_G16_mul2_G256_inv0 ^ z1911_assgn1911);
    assign z4705_assgn4705 = d0_G4_mul0_G16_mul2_G256_inv0;
    assign p1_domand2_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z1913_assgn1913);
    assign z4709_assgn4709 = d1_G4_mul0_G16_mul2_G256_inv0;
    assign p4_domand2_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z1915_assgn1915);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (i1_domand2_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_domand2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (i2_domand2_G4_mul0_G16_mul2_G256_inv0_reg ^ p4_domand2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z4721_assgn4721 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << z1925_assgn1925);
    assign z4725_assgn4725 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << z1927_assgn1927);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign z4733_assgn4733 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z1933_assgn1933);
    assign z4737_assgn4737 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z1935_assgn1935);
    assign z4741_assgn4741 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> z1937_assgn1937);
    assign z4745_assgn4745 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> z1939_assgn1939);
    assign z4749_assgn4749 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z1941_assgn1941);
    assign z4753_assgn4753 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z1943_assgn1943);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z4765_assgn4765 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << z1953_assgn1953);
    assign z4769_assgn4769 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << z1955_assgn1955);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign z4783_assgn4783 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z1967_assgn1967);
    assign z4787_assgn4787 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z1969_assgn1969);
    assign z4791_assgn4791 = dec_1_inp;
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> z1971_assgn1971);
    assign z4795_assgn4795 = dec_1_inp;
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> z1973_assgn1973);
    assign z4799_assgn4799 = dec_1_inp;
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z1975_assgn1975);
    assign z4803_assgn4803 = dec_1_inp;
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z1977_assgn1977);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ d1_G4_mul1_G16_mul2_G256_inv0);
    assign z0_domand0_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4829_assgn4829 = cxord_1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_domand0_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2001_assgn2001);
    assign z4833_assgn4833 = z0_domand0_G4_mul1_G16_mul2_G256_inv0;
    assign i1_domand0_G4_mul1_G16_mul2_G256_inv0 = (p2_domand0_G4_mul1_G16_mul2_G256_inv0 ^ z2003_assgn2003);
    assign z4837_assgn4837 = cxord_0_G4_mul1_G16_mul2_G256_inv0;
    assign p3_domand0_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2005_assgn2005);
    assign z4841_assgn4841 = z0_domand0_G4_mul1_G16_mul2_G256_inv0;
    assign i2_domand0_G4_mul1_G16_mul2_G256_inv0 = (p3_domand0_G4_mul1_G16_mul2_G256_inv0 ^ z2007_assgn2007);
    assign z4845_assgn4845 = cxord_0_G4_mul1_G16_mul2_G256_inv0;
    assign p1_domand0_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2009_assgn2009);
    assign z4849_assgn4849 = cxord_1_G4_mul1_G16_mul2_G256_inv0;
    assign p4_domand0_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2011_assgn2011);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (i1_domand0_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_domand0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (i2_domand0_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_domand0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z0_domand1_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4859_assgn4859 = c1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_domand1_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2019_assgn2019);
    assign z4863_assgn4863 = z0_domand1_G4_mul1_G16_mul2_G256_inv0;
    assign i1_domand1_G4_mul1_G16_mul2_G256_inv0 = (p2_domand1_G4_mul1_G16_mul2_G256_inv0 ^ z2021_assgn2021);
    assign z4867_assgn4867 = c0_G4_mul1_G16_mul2_G256_inv0;
    assign p3_domand1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2023_assgn2023);
    assign z4871_assgn4871 = z0_domand1_G4_mul1_G16_mul2_G256_inv0;
    assign i2_domand1_G4_mul1_G16_mul2_G256_inv0 = (p3_domand1_G4_mul1_G16_mul2_G256_inv0 ^ z2025_assgn2025);
    assign z4875_assgn4875 = c0_G4_mul1_G16_mul2_G256_inv0;
    assign p1_domand1_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2027_assgn2027);
    assign z4879_assgn4879 = c1_G4_mul1_G16_mul2_G256_inv0;
    assign p4_domand1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2029_assgn2029);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (i1_domand1_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_domand1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (i2_domand1_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_domand1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z0_domand2_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4893_assgn4893 = d1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_domand2_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2041_assgn2041);
    assign z4897_assgn4897 = z0_domand2_G4_mul1_G16_mul2_G256_inv0;
    assign i1_domand2_G4_mul1_G16_mul2_G256_inv0 = (p2_domand2_G4_mul1_G16_mul2_G256_inv0 ^ z2043_assgn2043);
    assign z4901_assgn4901 = d0_G4_mul1_G16_mul2_G256_inv0;
    assign p3_domand2_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2045_assgn2045);
    assign z4905_assgn4905 = z0_domand2_G4_mul1_G16_mul2_G256_inv0;
    assign i2_domand2_G4_mul1_G16_mul2_G256_inv0 = (p3_domand2_G4_mul1_G16_mul2_G256_inv0 ^ z2047_assgn2047);
    assign z4909_assgn4909 = d0_G4_mul1_G16_mul2_G256_inv0;
    assign p1_domand2_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2049_assgn2049);
    assign z4913_assgn4913 = d1_G4_mul1_G16_mul2_G256_inv0;
    assign p4_domand2_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2051_assgn2051);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (i1_domand2_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_domand2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (i2_domand2_G4_mul1_G16_mul2_G256_inv0_reg ^ p4_domand2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z4925_assgn4925 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << z2061_assgn2061);
    assign z4929_assgn4929 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << z2063_assgn2063);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r60_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r70_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r80_G16_mul2_G256_inv0 % dec_4_inp);
    assign z4947_assgn4947 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2079_assgn2079);
    assign z4951_assgn4951 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2081_assgn2081);
    assign z4955_assgn4955 = dec_1_inp;
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> z2083_assgn2083);
    assign z4959_assgn4959 = dec_1_inp;
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> z2085_assgn2085);
    assign z4963_assgn4963 = dec_1_inp;
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2087_assgn2087);
    assign z4967_assgn4967 = dec_1_inp;
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2089_assgn2089);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ d1_G4_mul2_G16_mul2_G256_inv0);
    assign z0_domand0_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign z4993_assgn4993 = cxord_1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_domand0_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2113_assgn2113);
    assign z4997_assgn4997 = z0_domand0_G4_mul2_G16_mul2_G256_inv0;
    assign i1_domand0_G4_mul2_G16_mul2_G256_inv0 = (p2_domand0_G4_mul2_G16_mul2_G256_inv0 ^ z2115_assgn2115);
    assign z5001_assgn5001 = cxord_0_G4_mul2_G16_mul2_G256_inv0;
    assign p3_domand0_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2117_assgn2117);
    assign z5005_assgn5005 = z0_domand0_G4_mul2_G16_mul2_G256_inv0;
    assign i2_domand0_G4_mul2_G16_mul2_G256_inv0 = (p3_domand0_G4_mul2_G16_mul2_G256_inv0 ^ z2119_assgn2119);
    assign z5009_assgn5009 = cxord_0_G4_mul2_G16_mul2_G256_inv0;
    assign p1_domand0_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2121_assgn2121);
    assign z5013_assgn5013 = cxord_1_G4_mul2_G16_mul2_G256_inv0;
    assign p4_domand0_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2123_assgn2123);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (i1_domand0_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_domand0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (i2_domand0_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_domand0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z0_domand1_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign z5023_assgn5023 = c1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_domand1_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2131_assgn2131);
    assign z5027_assgn5027 = z0_domand1_G4_mul2_G16_mul2_G256_inv0;
    assign i1_domand1_G4_mul2_G16_mul2_G256_inv0 = (p2_domand1_G4_mul2_G16_mul2_G256_inv0 ^ z2133_assgn2133);
    assign z5031_assgn5031 = c0_G4_mul2_G16_mul2_G256_inv0;
    assign p3_domand1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2135_assgn2135);
    assign z5035_assgn5035 = z0_domand1_G4_mul2_G16_mul2_G256_inv0;
    assign i2_domand1_G4_mul2_G16_mul2_G256_inv0 = (p3_domand1_G4_mul2_G16_mul2_G256_inv0 ^ z2137_assgn2137);
    assign z5039_assgn5039 = c0_G4_mul2_G16_mul2_G256_inv0;
    assign p1_domand1_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2139_assgn2139);
    assign z5043_assgn5043 = c1_G4_mul2_G16_mul2_G256_inv0;
    assign p4_domand1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2141_assgn2141);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (i1_domand1_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_domand1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (i2_domand1_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_domand1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z0_domand2_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign z5057_assgn5057 = d1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_domand2_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2153_assgn2153);
    assign z5061_assgn5061 = z0_domand2_G4_mul2_G16_mul2_G256_inv0;
    assign i1_domand2_G4_mul2_G16_mul2_G256_inv0 = (p2_domand2_G4_mul2_G16_mul2_G256_inv0 ^ z2155_assgn2155);
    assign z5065_assgn5065 = d0_G4_mul2_G16_mul2_G256_inv0;
    assign p3_domand2_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2157_assgn2157);
    assign z5069_assgn5069 = z0_domand2_G4_mul2_G16_mul2_G256_inv0;
    assign i2_domand2_G4_mul2_G16_mul2_G256_inv0 = (p3_domand2_G4_mul2_G16_mul2_G256_inv0 ^ z2159_assgn2159);
    assign z5073_assgn5073 = d0_G4_mul2_G16_mul2_G256_inv0;
    assign p1_domand2_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2161_assgn2161);
    assign z5077_assgn5077 = d1_G4_mul2_G16_mul2_G256_inv0;
    assign p4_domand2_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2163_assgn2163);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (i1_domand2_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_domand2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (i2_domand2_G4_mul2_G16_mul2_G256_inv0_reg ^ p4_domand2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z5089_assgn5089 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << z2173_assgn2173);
    assign z5093_assgn5093 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << z2175_assgn2175);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign z5105_assgn5105 = dec_2_inp;
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << z2185_assgn2185);
    assign z5109_assgn5109 = dec_2_inp;
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << z2187_assgn2187);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign z5117_assgn5117 = dec_4_inp;
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << z2193_assgn2193);
    assign z5121_assgn5121 = dec_4_inp;
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << z2195_assgn2195);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign z5133_assgn5133 = dec_1_inp;
    assign cond1_G256_newbasis1 = (t4 & z2205_assgn2205);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign z5141_assgn5141 = yxorb1_G256_newbasis1;
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * z2211_assgn2211);
    assign z5145_assgn5145 = tempy1_G256_newbasis1;
    assign tempybooloNegCond1_G256_newbasis1 = (z2214_assgn2214 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempybooloNegCond1_G256_newbasis1);
    assign z5151_assgn5151 = dec_1_inp;
    assign x1_G256_newbasis1 = (t4 >> z2217_assgn2217);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign z5157_assgn5157 = dec_1_inp;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & z2221_assgn2221);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign z5163_assgn5163 = dec_3_inp;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ z2225_assgn2225);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempybooloNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempybooloNegCond2_G256_newbasis1);
    assign z5173_assgn5173 = dec_1_inp;
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> z2233_assgn2233);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign z5179_assgn5179 = dec_1_inp;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & z2237_assgn2237);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign z5185_assgn5185 = dec_4_inp;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ z2241_assgn2241);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempybooloNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempybooloNegCond3_G256_newbasis1);
    assign z5195_assgn5195 = dec_1_inp;
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> z2249_assgn2249);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign z5201_assgn5201 = dec_1_inp;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & z2253_assgn2253);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign z5207_assgn5207 = dec_220_inp;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ z2257_assgn2257);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempybooloNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempybooloNegCond4_G256_newbasis1);
    assign z5217_assgn5217 = dec_1_inp;
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> z2265_assgn2265);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign z5223_assgn5223 = dec_1_inp;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & z2269_assgn2269);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign z5229_assgn5229 = dec_11_inp;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ z2273_assgn2273);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempybooloNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempybooloNegCond5_G256_newbasis1);
    assign z5239_assgn5239 = dec_1_inp;
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> z2281_assgn2281);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign z5245_assgn5245 = dec_1_inp;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & z2285_assgn2285);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign z5251_assgn5251 = dec_158_inp;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ z2289_assgn2289);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempybooloNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempybooloNegCond6_G256_newbasis1);
    assign z5261_assgn5261 = dec_1_inp;
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> z2297_assgn2297);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign z5267_assgn5267 = dec_1_inp;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & z2301_assgn2301);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign z5273_assgn5273 = dec_45_inp;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ z2305_assgn2305);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempybooloNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempybooloNegCond7_G256_newbasis1);
    assign z5283_assgn5283 = dec_1_inp;
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> z2313_assgn2313);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign z5289_assgn5289 = dec_1_inp;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & z2317_assgn2317);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign z5295_assgn5295 = dec_88_inp;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ z2321_assgn2321);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempybooloNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempybooloNegCond8_G256_newbasis1);
    assign z5305_assgn5305 = dec_1_inp;
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> z2329_assgn2329);
    assign t6 = y8_G256_newbasis1;
    assign z_y_G256_newbasis1 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z5315_assgn5315 = dec_1_inp;
    assign z_cond1_G256_newbasis1 = (t5 & z2337_assgn2337);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z5323_assgn5323 = z_yxorb1_G256_newbasis1;
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z2343_assgn2343);
    assign z5327_assgn5327 = z_tempy1_G256_newbasis1;
    assign z_tempybooloNegCond1_G256_newbasis1 = (z2346_assgn2346 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempybooloNegCond1_G256_newbasis1);
    assign z5333_assgn5333 = dec_1_inp;
    assign z_x1_G256_newbasis1 = (t5 >> z2349_assgn2349);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z5339_assgn5339 = dec_1_inp;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & z2353_assgn2353);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z5345_assgn5345 = dec_3_inp;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ z2357_assgn2357);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempybooloNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempybooloNegCond2_G256_newbasis1);
    assign z5355_assgn5355 = dec_1_inp;
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> z2365_assgn2365);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z5361_assgn5361 = dec_1_inp;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & z2369_assgn2369);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z5367_assgn5367 = dec_4_inp;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ z2373_assgn2373);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempybooloNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempybooloNegCond3_G256_newbasis1);
    assign z5377_assgn5377 = dec_1_inp;
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> z2381_assgn2381);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z5383_assgn5383 = dec_1_inp;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & z2385_assgn2385);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z5389_assgn5389 = dec_220_inp;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ z2389_assgn2389);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempybooloNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempybooloNegCond4_G256_newbasis1);
    assign z5399_assgn5399 = dec_1_inp;
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> z2397_assgn2397);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z5405_assgn5405 = dec_1_inp;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & z2401_assgn2401);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z5411_assgn5411 = dec_11_inp;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ z2405_assgn2405);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempybooloNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempybooloNegCond5_G256_newbasis1);
    assign z5421_assgn5421 = dec_1_inp;
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> z2413_assgn2413);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z5427_assgn5427 = dec_1_inp;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & z2417_assgn2417);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z5433_assgn5433 = dec_158_inp;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ z2421_assgn2421);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempybooloNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempybooloNegCond6_G256_newbasis1);
    assign z5443_assgn5443 = dec_1_inp;
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> z2429_assgn2429);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z5449_assgn5449 = dec_1_inp;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & z2433_assgn2433);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z5455_assgn5455 = dec_45_inp;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ z2437_assgn2437);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempybooloNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempybooloNegCond7_G256_newbasis1);
    assign z5465_assgn5465 = dec_1_inp;
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> z2445_assgn2445);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z5471_assgn5471 = dec_1_inp;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & z2449_assgn2449);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z5477_assgn5477 = dec_88_inp;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ z2453_assgn2453);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempybooloNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempybooloNegCond8_G256_newbasis1);
    assign z5487_assgn5487 = dec_1_inp;
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> z2461_assgn2461);
    assign t7 = z_y8_G256_newbasis1;
    assign z5493_assgn5493 = dec_99_inp;

    always @(posedge clk) begin
        z2721_assgn27210 <= z2721_assgn2721;
        z2721_assgn27211 <= z2721_assgn27210;
        z2721_assgn27212 <= z2721_assgn27211;
        x8_G256_newbasis0 <= z2721_assgn27212;
        z2853_assgn28530 <= z2853_assgn2853;
        z2853_assgn28531 <= z2853_assgn28530;
        z2853_assgn28532 <= z2853_assgn28531;
        z_x8_G256_newbasis0 <= z2853_assgn28532;
        i1_domand0_G4_mul0_G16_mul0_G256_inv0_reg <= i1_domand0_G4_mul0_G16_mul0_G256_inv0;
        p1_domand0_G4_mul0_G16_mul0_G256_inv0_reg <= p1_domand0_G4_mul0_G16_mul0_G256_inv0;
        i2_domand0_G4_mul0_G16_mul0_G256_inv0_reg <= i2_domand0_G4_mul0_G16_mul0_G256_inv0;
        p4_domand0_G4_mul0_G16_mul0_G256_inv0_reg <= p4_domand0_G4_mul0_G16_mul0_G256_inv0;
        i1_domand1_G4_mul0_G16_mul0_G256_inv0_reg <= i1_domand1_G4_mul0_G16_mul0_G256_inv0;
        p1_domand1_G4_mul0_G16_mul0_G256_inv0_reg <= p1_domand1_G4_mul0_G16_mul0_G256_inv0;
        i2_domand1_G4_mul0_G16_mul0_G256_inv0_reg <= i2_domand1_G4_mul0_G16_mul0_G256_inv0;
        p4_domand1_G4_mul0_G16_mul0_G256_inv0_reg <= p4_domand1_G4_mul0_G16_mul0_G256_inv0;
        i1_domand2_G4_mul0_G16_mul0_G256_inv0_reg <= i1_domand2_G4_mul0_G16_mul0_G256_inv0;
        p1_domand2_G4_mul0_G16_mul0_G256_inv0_reg <= p1_domand2_G4_mul0_G16_mul0_G256_inv0;
        i2_domand2_G4_mul0_G16_mul0_G256_inv0_reg <= i2_domand2_G4_mul0_G16_mul0_G256_inv0;
        p4_domand2_G4_mul0_G16_mul0_G256_inv0_reg <= p4_domand2_G4_mul0_G16_mul0_G256_inv0;
        dec_1_inp_reg <= dec_1_inp;
        dec_2_inp_reg <= dec_2_inp;
        i1_domand0_G4_mul1_G16_mul0_G256_inv0_reg <= i1_domand0_G4_mul1_G16_mul0_G256_inv0;
        p1_domand0_G4_mul1_G16_mul0_G256_inv0_reg <= p1_domand0_G4_mul1_G16_mul0_G256_inv0;
        i2_domand0_G4_mul1_G16_mul0_G256_inv0_reg <= i2_domand0_G4_mul1_G16_mul0_G256_inv0;
        p4_domand0_G4_mul1_G16_mul0_G256_inv0_reg <= p4_domand0_G4_mul1_G16_mul0_G256_inv0;
        i1_domand1_G4_mul1_G16_mul0_G256_inv0_reg <= i1_domand1_G4_mul1_G16_mul0_G256_inv0;
        p1_domand1_G4_mul1_G16_mul0_G256_inv0_reg <= p1_domand1_G4_mul1_G16_mul0_G256_inv0;
        i2_domand1_G4_mul1_G16_mul0_G256_inv0_reg <= i2_domand1_G4_mul1_G16_mul0_G256_inv0;
        p4_domand1_G4_mul1_G16_mul0_G256_inv0_reg <= p4_domand1_G4_mul1_G16_mul0_G256_inv0;
        i1_domand2_G4_mul1_G16_mul0_G256_inv0_reg <= i1_domand2_G4_mul1_G16_mul0_G256_inv0;
        p1_domand2_G4_mul1_G16_mul0_G256_inv0_reg <= p1_domand2_G4_mul1_G16_mul0_G256_inv0;
        i2_domand2_G4_mul1_G16_mul0_G256_inv0_reg <= i2_domand2_G4_mul1_G16_mul0_G256_inv0;
        p4_domand2_G4_mul1_G16_mul0_G256_inv0_reg <= p4_domand2_G4_mul1_G16_mul0_G256_inv0;
        i1_domand0_G4_mul2_G16_mul0_G256_inv0_reg <= i1_domand0_G4_mul2_G16_mul0_G256_inv0;
        p1_domand0_G4_mul2_G16_mul0_G256_inv0_reg <= p1_domand0_G4_mul2_G16_mul0_G256_inv0;
        i2_domand0_G4_mul2_G16_mul0_G256_inv0_reg <= i2_domand0_G4_mul2_G16_mul0_G256_inv0;
        p4_domand0_G4_mul2_G16_mul0_G256_inv0_reg <= p4_domand0_G4_mul2_G16_mul0_G256_inv0;
        i1_domand1_G4_mul2_G16_mul0_G256_inv0_reg <= i1_domand1_G4_mul2_G16_mul0_G256_inv0;
        p1_domand1_G4_mul2_G16_mul0_G256_inv0_reg <= p1_domand1_G4_mul2_G16_mul0_G256_inv0;
        i2_domand1_G4_mul2_G16_mul0_G256_inv0_reg <= i2_domand1_G4_mul2_G16_mul0_G256_inv0;
        p4_domand1_G4_mul2_G16_mul0_G256_inv0_reg <= p4_domand1_G4_mul2_G16_mul0_G256_inv0;
        i1_domand2_G4_mul2_G16_mul0_G256_inv0_reg <= i1_domand2_G4_mul2_G16_mul0_G256_inv0;
        p1_domand2_G4_mul2_G16_mul0_G256_inv0_reg <= p1_domand2_G4_mul2_G16_mul0_G256_inv0;
        i2_domand2_G4_mul2_G16_mul0_G256_inv0_reg <= i2_domand2_G4_mul2_G16_mul0_G256_inv0;
        p4_domand2_G4_mul2_G16_mul0_G256_inv0_reg <= p4_domand2_G4_mul2_G16_mul0_G256_inv0;
        c0_G256_inv0_reg <= c0_G256_inv0;
        c1_G256_inv0_reg <= c1_G256_inv0;
        dec_12_inp_reg <= dec_12_inp;
        dec_3_inp_reg <= dec_3_inp;
        z0_domand0_G4_mul3_G16_inv0_G256_inv0_reg <= z0_domand0_G4_mul3_G16_inv0_G256_inv0;
        i1_domand0_G4_mul3_G16_inv0_G256_inv0_reg <= i1_domand0_G4_mul3_G16_inv0_G256_inv0;
        p1_domand0_G4_mul3_G16_inv0_G256_inv0_reg <= p1_domand0_G4_mul3_G16_inv0_G256_inv0;
        i2_domand0_G4_mul3_G16_inv0_G256_inv0_reg <= i2_domand0_G4_mul3_G16_inv0_G256_inv0;
        p4_domand0_G4_mul3_G16_inv0_G256_inv0_reg <= p4_domand0_G4_mul3_G16_inv0_G256_inv0;
        z0_domand1_G4_mul3_G16_inv0_G256_inv0_reg <= z0_domand1_G4_mul3_G16_inv0_G256_inv0;
        i1_domand1_G4_mul3_G16_inv0_G256_inv0_reg <= i1_domand1_G4_mul3_G16_inv0_G256_inv0;
        p1_domand1_G4_mul3_G16_inv0_G256_inv0_reg <= p1_domand1_G4_mul3_G16_inv0_G256_inv0;
        i2_domand1_G4_mul3_G16_inv0_G256_inv0_reg <= i2_domand1_G4_mul3_G16_inv0_G256_inv0;
        p4_domand1_G4_mul3_G16_inv0_G256_inv0_reg <= p4_domand1_G4_mul3_G16_inv0_G256_inv0;
        z0_domand2_G4_mul3_G16_inv0_G256_inv0_reg <= z0_domand2_G4_mul3_G16_inv0_G256_inv0;
        i1_domand2_G4_mul3_G16_inv0_G256_inv0_reg <= i1_domand2_G4_mul3_G16_inv0_G256_inv0;
        p1_domand2_G4_mul3_G16_inv0_G256_inv0_reg <= p1_domand2_G4_mul3_G16_inv0_G256_inv0;
        i2_domand2_G4_mul3_G16_inv0_G256_inv0_reg <= i2_domand2_G4_mul3_G16_inv0_G256_inv0;
        p4_domand2_G4_mul3_G16_inv0_G256_inv0_reg <= p4_domand2_G4_mul3_G16_inv0_G256_inv0;
        z3569_assgn35690 <= z3569_assgn3569;
        z1101_assgn1101 <= z3569_assgn35690;
        z3573_assgn35730 <= z3573_assgn3573;
        z1103_assgn1103 <= z3573_assgn35730;
        c0_G16_inv0_G256_inv0_reg <= c0_G16_inv0_G256_inv0;
        c1_G16_inv0_G256_inv0_reg <= c1_G16_inv0_G256_inv0;
        z3585_assgn35850 <= z3585_assgn3585;
        z1113_assgn1113 <= z3585_assgn35850;
        z3589_assgn35890 <= z3589_assgn3589;
        z1115_assgn1115 <= z3589_assgn35890;
        z3593_assgn35930 <= z3593_assgn3593;
        z1117_assgn1117 <= z3593_assgn35930;
        z3597_assgn35970 <= z3597_assgn3597;
        z1119_assgn1119 <= z3597_assgn35970;
        z3601_assgn36010 <= z3601_assgn3601;
        z1121_assgn1121 <= z3601_assgn36010;
        z3605_assgn36050 <= z3605_assgn3605;
        z1123_assgn1123 <= z3605_assgn36050;
        z3609_assgn36090 <= z3609_assgn3609;
        z1125_assgn1125 <= z3609_assgn36090;
        z3613_assgn36130 <= z3613_assgn3613;
        z1127_assgn1127 <= z3613_assgn36130;
        z3627_assgn36270 <= z3627_assgn3627;
        z1139_assgn1139 <= z3627_assgn36270;
        z3631_assgn36310 <= z3631_assgn3631;
        z1141_assgn1141 <= z3631_assgn36310;
        z3635_assgn36350 <= z3635_assgn3635;
        z1143_assgn1143 <= z3635_assgn36350;
        z3639_assgn36390 <= z3639_assgn3639;
        z1145_assgn1145 <= z3639_assgn36390;
        z3643_assgn36430 <= z3643_assgn3643;
        z1147_assgn1147 <= z3643_assgn36430;
        z3647_assgn36470 <= z3647_assgn3647;
        z1149_assgn1149 <= z3647_assgn36470;
        cxord_1_G4_mul4_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul4_G16_inv0_G256_inv0;
        z3675_assgn36750 <= z3675_assgn3675;
        z1175_assgn1175 <= z3675_assgn36750;
        cxord_0_G4_mul4_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul4_G16_inv0_G256_inv0;
        z3681_assgn36810 <= z3681_assgn3681;
        z1179_assgn1179 <= z3681_assgn36810;
        i1_domand0_G4_mul4_G16_inv0_G256_inv0_reg <= i1_domand0_G4_mul4_G16_inv0_G256_inv0;
        p1_domand0_G4_mul4_G16_inv0_G256_inv0_reg <= p1_domand0_G4_mul4_G16_inv0_G256_inv0;
        i2_domand0_G4_mul4_G16_inv0_G256_inv0_reg <= i2_domand0_G4_mul4_G16_inv0_G256_inv0;
        p4_domand0_G4_mul4_G16_inv0_G256_inv0_reg <= p4_domand0_G4_mul4_G16_inv0_G256_inv0;
        c1_G4_mul4_G16_inv0_G256_inv0_reg <= c1_G4_mul4_G16_inv0_G256_inv0;
        z3697_assgn36970 <= z3697_assgn3697;
        z1193_assgn1193 <= z3697_assgn36970;
        c0_G4_mul4_G16_inv0_G256_inv0_reg <= c0_G4_mul4_G16_inv0_G256_inv0;
        z3703_assgn37030 <= z3703_assgn3703;
        z1197_assgn1197 <= z3703_assgn37030;
        i1_domand1_G4_mul4_G16_inv0_G256_inv0_reg <= i1_domand1_G4_mul4_G16_inv0_G256_inv0;
        p1_domand1_G4_mul4_G16_inv0_G256_inv0_reg <= p1_domand1_G4_mul4_G16_inv0_G256_inv0;
        i2_domand1_G4_mul4_G16_inv0_G256_inv0_reg <= i2_domand1_G4_mul4_G16_inv0_G256_inv0;
        p4_domand1_G4_mul4_G16_inv0_G256_inv0_reg <= p4_domand1_G4_mul4_G16_inv0_G256_inv0;
        d1_G4_mul4_G16_inv0_G256_inv0_reg <= d1_G4_mul4_G16_inv0_G256_inv0;
        z3723_assgn37230 <= z3723_assgn3723;
        z1215_assgn1215 <= z3723_assgn37230;
        d0_G4_mul4_G16_inv0_G256_inv0_reg <= d0_G4_mul4_G16_inv0_G256_inv0;
        z3729_assgn37290 <= z3729_assgn3729;
        z1219_assgn1219 <= z3729_assgn37290;
        i1_domand2_G4_mul4_G16_inv0_G256_inv0_reg <= i1_domand2_G4_mul4_G16_inv0_G256_inv0;
        p1_domand2_G4_mul4_G16_inv0_G256_inv0_reg <= p1_domand2_G4_mul4_G16_inv0_G256_inv0;
        i2_domand2_G4_mul4_G16_inv0_G256_inv0_reg <= i2_domand2_G4_mul4_G16_inv0_G256_inv0;
        p4_domand2_G4_mul4_G16_inv0_G256_inv0_reg <= p4_domand2_G4_mul4_G16_inv0_G256_inv0;
        z3745_assgn37450 <= z3745_assgn3745;
        z3745_assgn37451 <= z3745_assgn37450;
        z1233_assgn1233 <= z3745_assgn37451;
        z3749_assgn37490 <= z3749_assgn3749;
        z3749_assgn37491 <= z3749_assgn37490;
        z1235_assgn1235 <= z3749_assgn37491;
        z3763_assgn37630 <= z3763_assgn3763;
        z1247_assgn1247 <= z3763_assgn37630;
        z3767_assgn37670 <= z3767_assgn3767;
        z1249_assgn1249 <= z3767_assgn37670;
        z3771_assgn37710 <= z3771_assgn3771;
        z1251_assgn1251 <= z3771_assgn37710;
        z3775_assgn37750 <= z3775_assgn3775;
        z1253_assgn1253 <= z3775_assgn37750;
        z3779_assgn37790 <= z3779_assgn3779;
        z1255_assgn1255 <= z3779_assgn37790;
        z3783_assgn37830 <= z3783_assgn3783;
        z1257_assgn1257 <= z3783_assgn37830;
        cxord_1_G4_mul5_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul5_G16_inv0_G256_inv0;
        z3811_assgn38110 <= z3811_assgn3811;
        z1283_assgn1283 <= z3811_assgn38110;
        cxord_0_G4_mul5_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul5_G16_inv0_G256_inv0;
        z3817_assgn38170 <= z3817_assgn3817;
        z1287_assgn1287 <= z3817_assgn38170;
        i1_domand0_G4_mul5_G16_inv0_G256_inv0_reg <= i1_domand0_G4_mul5_G16_inv0_G256_inv0;
        p1_domand0_G4_mul5_G16_inv0_G256_inv0_reg <= p1_domand0_G4_mul5_G16_inv0_G256_inv0;
        i2_domand0_G4_mul5_G16_inv0_G256_inv0_reg <= i2_domand0_G4_mul5_G16_inv0_G256_inv0;
        p4_domand0_G4_mul5_G16_inv0_G256_inv0_reg <= p4_domand0_G4_mul5_G16_inv0_G256_inv0;
        c1_G4_mul5_G16_inv0_G256_inv0_reg <= c1_G4_mul5_G16_inv0_G256_inv0;
        z3833_assgn38330 <= z3833_assgn3833;
        z1301_assgn1301 <= z3833_assgn38330;
        c0_G4_mul5_G16_inv0_G256_inv0_reg <= c0_G4_mul5_G16_inv0_G256_inv0;
        z3839_assgn38390 <= z3839_assgn3839;
        z1305_assgn1305 <= z3839_assgn38390;
        i1_domand1_G4_mul5_G16_inv0_G256_inv0_reg <= i1_domand1_G4_mul5_G16_inv0_G256_inv0;
        p1_domand1_G4_mul5_G16_inv0_G256_inv0_reg <= p1_domand1_G4_mul5_G16_inv0_G256_inv0;
        i2_domand1_G4_mul5_G16_inv0_G256_inv0_reg <= i2_domand1_G4_mul5_G16_inv0_G256_inv0;
        p4_domand1_G4_mul5_G16_inv0_G256_inv0_reg <= p4_domand1_G4_mul5_G16_inv0_G256_inv0;
        d1_G4_mul5_G16_inv0_G256_inv0_reg <= d1_G4_mul5_G16_inv0_G256_inv0;
        z3859_assgn38590 <= z3859_assgn3859;
        z1323_assgn1323 <= z3859_assgn38590;
        d0_G4_mul5_G16_inv0_G256_inv0_reg <= d0_G4_mul5_G16_inv0_G256_inv0;
        z3865_assgn38650 <= z3865_assgn3865;
        z1327_assgn1327 <= z3865_assgn38650;
        i1_domand2_G4_mul5_G16_inv0_G256_inv0_reg <= i1_domand2_G4_mul5_G16_inv0_G256_inv0;
        p1_domand2_G4_mul5_G16_inv0_G256_inv0_reg <= p1_domand2_G4_mul5_G16_inv0_G256_inv0;
        i2_domand2_G4_mul5_G16_inv0_G256_inv0_reg <= i2_domand2_G4_mul5_G16_inv0_G256_inv0;
        p4_domand2_G4_mul5_G16_inv0_G256_inv0_reg <= p4_domand2_G4_mul5_G16_inv0_G256_inv0;
        z3881_assgn38810 <= z3881_assgn3881;
        z3881_assgn38811 <= z3881_assgn38810;
        z1341_assgn1341 <= z3881_assgn38811;
        z3885_assgn38850 <= z3885_assgn3885;
        z3885_assgn38851 <= z3885_assgn38850;
        z1343_assgn1343 <= z3885_assgn38851;
        z3893_assgn38930 <= z3893_assgn3893;
        z3893_assgn38931 <= z3893_assgn38930;
        z1349_assgn1349 <= z3893_assgn38931;
        z3897_assgn38970 <= z3897_assgn3897;
        z3897_assgn38971 <= z3897_assgn38970;
        z1351_assgn1351 <= z3897_assgn38971;
        z3923_assgn39230 <= z3923_assgn3923;
        z3923_assgn39231 <= z3923_assgn39230;
        z1375_assgn1375 <= z3923_assgn39231;
        z3927_assgn39270 <= z3927_assgn3927;
        z3927_assgn39271 <= z3927_assgn39270;
        z1377_assgn1377 <= z3927_assgn39271;
        z3931_assgn39310 <= z3931_assgn3931;
        z3931_assgn39311 <= z3931_assgn39310;
        z1379_assgn1379 <= z3931_assgn39311;
        z3935_assgn39350 <= z3935_assgn3935;
        z3935_assgn39351 <= z3935_assgn39350;
        z1381_assgn1381 <= z3935_assgn39351;
        z3939_assgn39390 <= z3939_assgn3939;
        z3939_assgn39391 <= z3939_assgn39390;
        z1383_assgn1383 <= z3939_assgn39391;
        z3943_assgn39430 <= z3943_assgn3943;
        z3943_assgn39431 <= z3943_assgn39430;
        z1385_assgn1385 <= z3943_assgn39431;
        z3973_assgn39730 <= z3973_assgn3973;
        z3973_assgn39731 <= z3973_assgn39730;
        z1413_assgn1413 <= z3973_assgn39731;
        z3977_assgn39770 <= z3977_assgn3977;
        z3977_assgn39771 <= z3977_assgn39770;
        z1415_assgn1415 <= z3977_assgn39771;
        z3981_assgn39810 <= z3981_assgn3981;
        z3981_assgn39811 <= z3981_assgn39810;
        z1417_assgn1417 <= z3981_assgn39811;
        z3985_assgn39850 <= z3985_assgn3985;
        z3985_assgn39851 <= z3985_assgn39850;
        z1419_assgn1419 <= z3985_assgn39851;
        z3989_assgn39890 <= z3989_assgn3989;
        z3989_assgn39891 <= z3989_assgn39890;
        z1421_assgn1421 <= z3989_assgn39891;
        z3993_assgn39930 <= z3993_assgn3993;
        z3993_assgn39931 <= z3993_assgn39930;
        z1423_assgn1423 <= z3993_assgn39931;
        z4019_assgn40190 <= z4019_assgn4019;
        z4019_assgn40191 <= z4019_assgn40190;
        z1447_assgn1447 <= z4019_assgn40191;
        z4023_assgn40230 <= z4023_assgn4023;
        z4023_assgn40231 <= z4023_assgn40230;
        z1449_assgn1449 <= z4023_assgn40231;
        z4027_assgn40270 <= z4027_assgn4027;
        z4027_assgn40271 <= z4027_assgn40270;
        z1451_assgn1451 <= z4027_assgn40271;
        z4031_assgn40310 <= z4031_assgn4031;
        z4031_assgn40311 <= z4031_assgn40310;
        z1453_assgn1453 <= z4031_assgn40311;
        z4035_assgn40350 <= z4035_assgn4035;
        z4035_assgn40351 <= z4035_assgn40350;
        z1455_assgn1455 <= z4035_assgn40351;
        z4039_assgn40390 <= z4039_assgn4039;
        z4039_assgn40391 <= z4039_assgn40390;
        z1457_assgn1457 <= z4039_assgn40391;
        i1_domand0_G4_mul0_G16_mul1_G256_inv0_reg <= i1_domand0_G4_mul0_G16_mul1_G256_inv0;
        p1_domand0_G4_mul0_G16_mul1_G256_inv0_reg <= p1_domand0_G4_mul0_G16_mul1_G256_inv0;
        i2_domand0_G4_mul0_G16_mul1_G256_inv0_reg <= i2_domand0_G4_mul0_G16_mul1_G256_inv0;
        p4_domand0_G4_mul0_G16_mul1_G256_inv0_reg <= p4_domand0_G4_mul0_G16_mul1_G256_inv0;
        z4049_assgn40490 <= z4049_assgn4049;
        z4049_assgn40491 <= z4049_assgn40490;
        z1465_assgn1465 <= z4049_assgn40491;
        z4053_assgn40530 <= z4053_assgn4053;
        z4053_assgn40531 <= z4053_assgn40530;
        z1467_assgn1467 <= z4053_assgn40531;
        z4057_assgn40570 <= z4057_assgn4057;
        z4057_assgn40571 <= z4057_assgn40570;
        z1469_assgn1469 <= z4057_assgn40571;
        z4061_assgn40610 <= z4061_assgn4061;
        z4061_assgn40611 <= z4061_assgn40610;
        z1471_assgn1471 <= z4061_assgn40611;
        z4065_assgn40650 <= z4065_assgn4065;
        z4065_assgn40651 <= z4065_assgn40650;
        z1473_assgn1473 <= z4065_assgn40651;
        z4069_assgn40690 <= z4069_assgn4069;
        z4069_assgn40691 <= z4069_assgn40690;
        z1475_assgn1475 <= z4069_assgn40691;
        i1_domand1_G4_mul0_G16_mul1_G256_inv0_reg <= i1_domand1_G4_mul0_G16_mul1_G256_inv0;
        p1_domand1_G4_mul0_G16_mul1_G256_inv0_reg <= p1_domand1_G4_mul0_G16_mul1_G256_inv0;
        i2_domand1_G4_mul0_G16_mul1_G256_inv0_reg <= i2_domand1_G4_mul0_G16_mul1_G256_inv0;
        p4_domand1_G4_mul0_G16_mul1_G256_inv0_reg <= p4_domand1_G4_mul0_G16_mul1_G256_inv0;
        z4083_assgn40830 <= z4083_assgn4083;
        z4083_assgn40831 <= z4083_assgn40830;
        z1487_assgn1487 <= z4083_assgn40831;
        z4087_assgn40870 <= z4087_assgn4087;
        z4087_assgn40871 <= z4087_assgn40870;
        z1489_assgn1489 <= z4087_assgn40871;
        z4091_assgn40910 <= z4091_assgn4091;
        z4091_assgn40911 <= z4091_assgn40910;
        z1491_assgn1491 <= z4091_assgn40911;
        z4095_assgn40950 <= z4095_assgn4095;
        z4095_assgn40951 <= z4095_assgn40950;
        z1493_assgn1493 <= z4095_assgn40951;
        z4099_assgn40990 <= z4099_assgn4099;
        z4099_assgn40991 <= z4099_assgn40990;
        z1495_assgn1495 <= z4099_assgn40991;
        z4103_assgn41030 <= z4103_assgn4103;
        z4103_assgn41031 <= z4103_assgn41030;
        z1497_assgn1497 <= z4103_assgn41031;
        i1_domand2_G4_mul0_G16_mul1_G256_inv0_reg <= i1_domand2_G4_mul0_G16_mul1_G256_inv0;
        p1_domand2_G4_mul0_G16_mul1_G256_inv0_reg <= p1_domand2_G4_mul0_G16_mul1_G256_inv0;
        i2_domand2_G4_mul0_G16_mul1_G256_inv0_reg <= i2_domand2_G4_mul0_G16_mul1_G256_inv0;
        p4_domand2_G4_mul0_G16_mul1_G256_inv0_reg <= p4_domand2_G4_mul0_G16_mul1_G256_inv0;
        z4115_assgn41150 <= z4115_assgn4115;
        z4115_assgn41151 <= z4115_assgn41150;
        z4115_assgn41152 <= z4115_assgn41151;
        z1507_assgn1507 <= z4115_assgn41152;
        z4119_assgn41190 <= z4119_assgn4119;
        z4119_assgn41191 <= z4119_assgn41190;
        z4119_assgn41192 <= z4119_assgn41191;
        z1509_assgn1509 <= z4119_assgn41192;
        z4127_assgn41270 <= z4127_assgn4127;
        z4127_assgn41271 <= z4127_assgn41270;
        z4127_assgn41272 <= z4127_assgn41271;
        z1515_assgn1515 <= z4127_assgn41272;
        z4131_assgn41310 <= z4131_assgn4131;
        z4131_assgn41311 <= z4131_assgn41310;
        z4131_assgn41312 <= z4131_assgn41311;
        z1517_assgn1517 <= z4131_assgn41312;
        z4135_assgn41350 <= z4135_assgn4135;
        z4135_assgn41351 <= z4135_assgn41350;
        z4135_assgn41352 <= z4135_assgn41351;
        z1519_assgn1519 <= z4135_assgn41352;
        z4139_assgn41390 <= z4139_assgn4139;
        z4139_assgn41391 <= z4139_assgn41390;
        z4139_assgn41392 <= z4139_assgn41391;
        z1521_assgn1521 <= z4139_assgn41392;
        z4143_assgn41430 <= z4143_assgn4143;
        z4143_assgn41431 <= z4143_assgn41430;
        z4143_assgn41432 <= z4143_assgn41431;
        z1523_assgn1523 <= z4143_assgn41432;
        z4147_assgn41470 <= z4147_assgn4147;
        z4147_assgn41471 <= z4147_assgn41470;
        z4147_assgn41472 <= z4147_assgn41471;
        z1525_assgn1525 <= z4147_assgn41472;
        z4159_assgn41590 <= z4159_assgn4159;
        z4159_assgn41591 <= z4159_assgn41590;
        z4159_assgn41592 <= z4159_assgn41591;
        z1535_assgn1535 <= z4159_assgn41592;
        z4163_assgn41630 <= z4163_assgn4163;
        z4163_assgn41631 <= z4163_assgn41630;
        z4163_assgn41632 <= z4163_assgn41631;
        z1537_assgn1537 <= z4163_assgn41632;
        z4177_assgn41770 <= z4177_assgn4177;
        z4177_assgn41771 <= z4177_assgn41770;
        z1549_assgn1549 <= z4177_assgn41771;
        z4181_assgn41810 <= z4181_assgn4181;
        z4181_assgn41811 <= z4181_assgn41810;
        z1551_assgn1551 <= z4181_assgn41811;
        z4185_assgn41850 <= z4185_assgn4185;
        z4185_assgn41851 <= z4185_assgn41850;
        z1553_assgn1553 <= z4185_assgn41851;
        z4189_assgn41890 <= z4189_assgn4189;
        z4189_assgn41891 <= z4189_assgn41890;
        z1555_assgn1555 <= z4189_assgn41891;
        z4193_assgn41930 <= z4193_assgn4193;
        z4193_assgn41931 <= z4193_assgn41930;
        z1557_assgn1557 <= z4193_assgn41931;
        z4197_assgn41970 <= z4197_assgn4197;
        z4197_assgn41971 <= z4197_assgn41970;
        z1559_assgn1559 <= z4197_assgn41971;
        z4223_assgn42230 <= z4223_assgn4223;
        z4223_assgn42231 <= z4223_assgn42230;
        z1583_assgn1583 <= z4223_assgn42231;
        z4227_assgn42270 <= z4227_assgn4227;
        z4227_assgn42271 <= z4227_assgn42270;
        z1585_assgn1585 <= z4227_assgn42271;
        z4231_assgn42310 <= z4231_assgn4231;
        z4231_assgn42311 <= z4231_assgn42310;
        z1587_assgn1587 <= z4231_assgn42311;
        z4235_assgn42350 <= z4235_assgn4235;
        z4235_assgn42351 <= z4235_assgn42350;
        z1589_assgn1589 <= z4235_assgn42351;
        z4239_assgn42390 <= z4239_assgn4239;
        z4239_assgn42391 <= z4239_assgn42390;
        z1591_assgn1591 <= z4239_assgn42391;
        z4243_assgn42430 <= z4243_assgn4243;
        z4243_assgn42431 <= z4243_assgn42430;
        z1593_assgn1593 <= z4243_assgn42431;
        i1_domand0_G4_mul1_G16_mul1_G256_inv0_reg <= i1_domand0_G4_mul1_G16_mul1_G256_inv0;
        p1_domand0_G4_mul1_G16_mul1_G256_inv0_reg <= p1_domand0_G4_mul1_G16_mul1_G256_inv0;
        i2_domand0_G4_mul1_G16_mul1_G256_inv0_reg <= i2_domand0_G4_mul1_G16_mul1_G256_inv0;
        p4_domand0_G4_mul1_G16_mul1_G256_inv0_reg <= p4_domand0_G4_mul1_G16_mul1_G256_inv0;
        z4253_assgn42530 <= z4253_assgn4253;
        z4253_assgn42531 <= z4253_assgn42530;
        z1601_assgn1601 <= z4253_assgn42531;
        z4257_assgn42570 <= z4257_assgn4257;
        z4257_assgn42571 <= z4257_assgn42570;
        z1603_assgn1603 <= z4257_assgn42571;
        z4261_assgn42610 <= z4261_assgn4261;
        z4261_assgn42611 <= z4261_assgn42610;
        z1605_assgn1605 <= z4261_assgn42611;
        z4265_assgn42650 <= z4265_assgn4265;
        z4265_assgn42651 <= z4265_assgn42650;
        z1607_assgn1607 <= z4265_assgn42651;
        z4269_assgn42690 <= z4269_assgn4269;
        z4269_assgn42691 <= z4269_assgn42690;
        z1609_assgn1609 <= z4269_assgn42691;
        z4273_assgn42730 <= z4273_assgn4273;
        z4273_assgn42731 <= z4273_assgn42730;
        z1611_assgn1611 <= z4273_assgn42731;
        i1_domand1_G4_mul1_G16_mul1_G256_inv0_reg <= i1_domand1_G4_mul1_G16_mul1_G256_inv0;
        p1_domand1_G4_mul1_G16_mul1_G256_inv0_reg <= p1_domand1_G4_mul1_G16_mul1_G256_inv0;
        i2_domand1_G4_mul1_G16_mul1_G256_inv0_reg <= i2_domand1_G4_mul1_G16_mul1_G256_inv0;
        p4_domand1_G4_mul1_G16_mul1_G256_inv0_reg <= p4_domand1_G4_mul1_G16_mul1_G256_inv0;
        z4287_assgn42870 <= z4287_assgn4287;
        z4287_assgn42871 <= z4287_assgn42870;
        z1623_assgn1623 <= z4287_assgn42871;
        z4291_assgn42910 <= z4291_assgn4291;
        z4291_assgn42911 <= z4291_assgn42910;
        z1625_assgn1625 <= z4291_assgn42911;
        z4295_assgn42950 <= z4295_assgn4295;
        z4295_assgn42951 <= z4295_assgn42950;
        z1627_assgn1627 <= z4295_assgn42951;
        z4299_assgn42990 <= z4299_assgn4299;
        z4299_assgn42991 <= z4299_assgn42990;
        z1629_assgn1629 <= z4299_assgn42991;
        z4303_assgn43030 <= z4303_assgn4303;
        z4303_assgn43031 <= z4303_assgn43030;
        z1631_assgn1631 <= z4303_assgn43031;
        z4307_assgn43070 <= z4307_assgn4307;
        z4307_assgn43071 <= z4307_assgn43070;
        z1633_assgn1633 <= z4307_assgn43071;
        i1_domand2_G4_mul1_G16_mul1_G256_inv0_reg <= i1_domand2_G4_mul1_G16_mul1_G256_inv0;
        p1_domand2_G4_mul1_G16_mul1_G256_inv0_reg <= p1_domand2_G4_mul1_G16_mul1_G256_inv0;
        i2_domand2_G4_mul1_G16_mul1_G256_inv0_reg <= i2_domand2_G4_mul1_G16_mul1_G256_inv0;
        p4_domand2_G4_mul1_G16_mul1_G256_inv0_reg <= p4_domand2_G4_mul1_G16_mul1_G256_inv0;
        z4319_assgn43190 <= z4319_assgn4319;
        z4319_assgn43191 <= z4319_assgn43190;
        z4319_assgn43192 <= z4319_assgn43191;
        z1643_assgn1643 <= z4319_assgn43192;
        z4323_assgn43230 <= z4323_assgn4323;
        z4323_assgn43231 <= z4323_assgn43230;
        z4323_assgn43232 <= z4323_assgn43231;
        z1645_assgn1645 <= z4323_assgn43232;
        z4341_assgn43410 <= z4341_assgn4341;
        z4341_assgn43411 <= z4341_assgn43410;
        z1661_assgn1661 <= z4341_assgn43411;
        z4345_assgn43450 <= z4345_assgn4345;
        z4345_assgn43451 <= z4345_assgn43450;
        z1663_assgn1663 <= z4345_assgn43451;
        z4349_assgn43490 <= z4349_assgn4349;
        z4349_assgn43491 <= z4349_assgn43490;
        z1665_assgn1665 <= z4349_assgn43491;
        z4353_assgn43530 <= z4353_assgn4353;
        z4353_assgn43531 <= z4353_assgn43530;
        z1667_assgn1667 <= z4353_assgn43531;
        z4357_assgn43570 <= z4357_assgn4357;
        z4357_assgn43571 <= z4357_assgn43570;
        z1669_assgn1669 <= z4357_assgn43571;
        z4361_assgn43610 <= z4361_assgn4361;
        z4361_assgn43611 <= z4361_assgn43610;
        z1671_assgn1671 <= z4361_assgn43611;
        z4387_assgn43870 <= z4387_assgn4387;
        z4387_assgn43871 <= z4387_assgn43870;
        z1695_assgn1695 <= z4387_assgn43871;
        z4391_assgn43910 <= z4391_assgn4391;
        z4391_assgn43911 <= z4391_assgn43910;
        z1697_assgn1697 <= z4391_assgn43911;
        z4395_assgn43950 <= z4395_assgn4395;
        z4395_assgn43951 <= z4395_assgn43950;
        z1699_assgn1699 <= z4395_assgn43951;
        z4399_assgn43990 <= z4399_assgn4399;
        z4399_assgn43991 <= z4399_assgn43990;
        z1701_assgn1701 <= z4399_assgn43991;
        z4403_assgn44030 <= z4403_assgn4403;
        z4403_assgn44031 <= z4403_assgn44030;
        z1703_assgn1703 <= z4403_assgn44031;
        z4407_assgn44070 <= z4407_assgn4407;
        z4407_assgn44071 <= z4407_assgn44070;
        z1705_assgn1705 <= z4407_assgn44071;
        i1_domand0_G4_mul2_G16_mul1_G256_inv0_reg <= i1_domand0_G4_mul2_G16_mul1_G256_inv0;
        p1_domand0_G4_mul2_G16_mul1_G256_inv0_reg <= p1_domand0_G4_mul2_G16_mul1_G256_inv0;
        i2_domand0_G4_mul2_G16_mul1_G256_inv0_reg <= i2_domand0_G4_mul2_G16_mul1_G256_inv0;
        p4_domand0_G4_mul2_G16_mul1_G256_inv0_reg <= p4_domand0_G4_mul2_G16_mul1_G256_inv0;
        z4417_assgn44170 <= z4417_assgn4417;
        z4417_assgn44171 <= z4417_assgn44170;
        z1713_assgn1713 <= z4417_assgn44171;
        z4421_assgn44210 <= z4421_assgn4421;
        z4421_assgn44211 <= z4421_assgn44210;
        z1715_assgn1715 <= z4421_assgn44211;
        z4425_assgn44250 <= z4425_assgn4425;
        z4425_assgn44251 <= z4425_assgn44250;
        z1717_assgn1717 <= z4425_assgn44251;
        z4429_assgn44290 <= z4429_assgn4429;
        z4429_assgn44291 <= z4429_assgn44290;
        z1719_assgn1719 <= z4429_assgn44291;
        z4433_assgn44330 <= z4433_assgn4433;
        z4433_assgn44331 <= z4433_assgn44330;
        z1721_assgn1721 <= z4433_assgn44331;
        z4437_assgn44370 <= z4437_assgn4437;
        z4437_assgn44371 <= z4437_assgn44370;
        z1723_assgn1723 <= z4437_assgn44371;
        i1_domand1_G4_mul2_G16_mul1_G256_inv0_reg <= i1_domand1_G4_mul2_G16_mul1_G256_inv0;
        p1_domand1_G4_mul2_G16_mul1_G256_inv0_reg <= p1_domand1_G4_mul2_G16_mul1_G256_inv0;
        i2_domand1_G4_mul2_G16_mul1_G256_inv0_reg <= i2_domand1_G4_mul2_G16_mul1_G256_inv0;
        p4_domand1_G4_mul2_G16_mul1_G256_inv0_reg <= p4_domand1_G4_mul2_G16_mul1_G256_inv0;
        z4451_assgn44510 <= z4451_assgn4451;
        z4451_assgn44511 <= z4451_assgn44510;
        z1735_assgn1735 <= z4451_assgn44511;
        z4455_assgn44550 <= z4455_assgn4455;
        z4455_assgn44551 <= z4455_assgn44550;
        z1737_assgn1737 <= z4455_assgn44551;
        z4459_assgn44590 <= z4459_assgn4459;
        z4459_assgn44591 <= z4459_assgn44590;
        z1739_assgn1739 <= z4459_assgn44591;
        z4463_assgn44630 <= z4463_assgn4463;
        z4463_assgn44631 <= z4463_assgn44630;
        z1741_assgn1741 <= z4463_assgn44631;
        z4467_assgn44670 <= z4467_assgn4467;
        z4467_assgn44671 <= z4467_assgn44670;
        z1743_assgn1743 <= z4467_assgn44671;
        z4471_assgn44710 <= z4471_assgn4471;
        z4471_assgn44711 <= z4471_assgn44710;
        z1745_assgn1745 <= z4471_assgn44711;
        i1_domand2_G4_mul2_G16_mul1_G256_inv0_reg <= i1_domand2_G4_mul2_G16_mul1_G256_inv0;
        p1_domand2_G4_mul2_G16_mul1_G256_inv0_reg <= p1_domand2_G4_mul2_G16_mul1_G256_inv0;
        i2_domand2_G4_mul2_G16_mul1_G256_inv0_reg <= i2_domand2_G4_mul2_G16_mul1_G256_inv0;
        p4_domand2_G4_mul2_G16_mul1_G256_inv0_reg <= p4_domand2_G4_mul2_G16_mul1_G256_inv0;
        z4483_assgn44830 <= z4483_assgn4483;
        z4483_assgn44831 <= z4483_assgn44830;
        z4483_assgn44832 <= z4483_assgn44831;
        z1755_assgn1755 <= z4483_assgn44832;
        z4487_assgn44870 <= z4487_assgn4487;
        z4487_assgn44871 <= z4487_assgn44870;
        z4487_assgn44872 <= z4487_assgn44871;
        z1757_assgn1757 <= z4487_assgn44872;
        z4499_assgn44990 <= z4499_assgn4499;
        z4499_assgn44991 <= z4499_assgn44990;
        z4499_assgn44992 <= z4499_assgn44991;
        z1767_assgn1767 <= z4499_assgn44992;
        z4503_assgn45030 <= z4503_assgn4503;
        z4503_assgn45031 <= z4503_assgn45030;
        z4503_assgn45032 <= z4503_assgn45031;
        z1769_assgn1769 <= z4503_assgn45032;
        z4529_assgn45290 <= z4529_assgn4529;
        z4529_assgn45291 <= z4529_assgn45290;
        z1793_assgn1793 <= z4529_assgn45291;
        z4533_assgn45330 <= z4533_assgn4533;
        z4533_assgn45331 <= z4533_assgn45330;
        z1795_assgn1795 <= z4533_assgn45331;
        z4537_assgn45370 <= z4537_assgn4537;
        z4537_assgn45371 <= z4537_assgn45370;
        z1797_assgn1797 <= z4537_assgn45371;
        z4541_assgn45410 <= z4541_assgn4541;
        z4541_assgn45411 <= z4541_assgn45410;
        z1799_assgn1799 <= z4541_assgn45411;
        z4545_assgn45450 <= z4545_assgn4545;
        z4545_assgn45451 <= z4545_assgn45450;
        z1801_assgn1801 <= z4545_assgn45451;
        z4549_assgn45490 <= z4549_assgn4549;
        z4549_assgn45491 <= z4549_assgn45490;
        z1803_assgn1803 <= z4549_assgn45491;
        z4579_assgn45790 <= z4579_assgn4579;
        z4579_assgn45791 <= z4579_assgn45790;
        z1831_assgn1831 <= z4579_assgn45791;
        z4583_assgn45830 <= z4583_assgn4583;
        z4583_assgn45831 <= z4583_assgn45830;
        z1833_assgn1833 <= z4583_assgn45831;
        z4587_assgn45870 <= z4587_assgn4587;
        z4587_assgn45871 <= z4587_assgn45870;
        z1835_assgn1835 <= z4587_assgn45871;
        z4591_assgn45910 <= z4591_assgn4591;
        z4591_assgn45911 <= z4591_assgn45910;
        z1837_assgn1837 <= z4591_assgn45911;
        z4595_assgn45950 <= z4595_assgn4595;
        z4595_assgn45951 <= z4595_assgn45950;
        z1839_assgn1839 <= z4595_assgn45951;
        z4599_assgn45990 <= z4599_assgn4599;
        z4599_assgn45991 <= z4599_assgn45990;
        z1841_assgn1841 <= z4599_assgn45991;
        z4625_assgn46250 <= z4625_assgn4625;
        z4625_assgn46251 <= z4625_assgn46250;
        z1865_assgn1865 <= z4625_assgn46251;
        z4629_assgn46290 <= z4629_assgn4629;
        z4629_assgn46291 <= z4629_assgn46290;
        z1867_assgn1867 <= z4629_assgn46291;
        z4633_assgn46330 <= z4633_assgn4633;
        z4633_assgn46331 <= z4633_assgn46330;
        z1869_assgn1869 <= z4633_assgn46331;
        z4637_assgn46370 <= z4637_assgn4637;
        z4637_assgn46371 <= z4637_assgn46370;
        z1871_assgn1871 <= z4637_assgn46371;
        z4641_assgn46410 <= z4641_assgn4641;
        z4641_assgn46411 <= z4641_assgn46410;
        z1873_assgn1873 <= z4641_assgn46411;
        z4645_assgn46450 <= z4645_assgn4645;
        z4645_assgn46451 <= z4645_assgn46450;
        z1875_assgn1875 <= z4645_assgn46451;
        i1_domand0_G4_mul0_G16_mul2_G256_inv0_reg <= i1_domand0_G4_mul0_G16_mul2_G256_inv0;
        p1_domand0_G4_mul0_G16_mul2_G256_inv0_reg <= p1_domand0_G4_mul0_G16_mul2_G256_inv0;
        i2_domand0_G4_mul0_G16_mul2_G256_inv0_reg <= i2_domand0_G4_mul0_G16_mul2_G256_inv0;
        p4_domand0_G4_mul0_G16_mul2_G256_inv0_reg <= p4_domand0_G4_mul0_G16_mul2_G256_inv0;
        z4655_assgn46550 <= z4655_assgn4655;
        z4655_assgn46551 <= z4655_assgn46550;
        z1883_assgn1883 <= z4655_assgn46551;
        z4659_assgn46590 <= z4659_assgn4659;
        z4659_assgn46591 <= z4659_assgn46590;
        z1885_assgn1885 <= z4659_assgn46591;
        z4663_assgn46630 <= z4663_assgn4663;
        z4663_assgn46631 <= z4663_assgn46630;
        z1887_assgn1887 <= z4663_assgn46631;
        z4667_assgn46670 <= z4667_assgn4667;
        z4667_assgn46671 <= z4667_assgn46670;
        z1889_assgn1889 <= z4667_assgn46671;
        z4671_assgn46710 <= z4671_assgn4671;
        z4671_assgn46711 <= z4671_assgn46710;
        z1891_assgn1891 <= z4671_assgn46711;
        z4675_assgn46750 <= z4675_assgn4675;
        z4675_assgn46751 <= z4675_assgn46750;
        z1893_assgn1893 <= z4675_assgn46751;
        i1_domand1_G4_mul0_G16_mul2_G256_inv0_reg <= i1_domand1_G4_mul0_G16_mul2_G256_inv0;
        p1_domand1_G4_mul0_G16_mul2_G256_inv0_reg <= p1_domand1_G4_mul0_G16_mul2_G256_inv0;
        i2_domand1_G4_mul0_G16_mul2_G256_inv0_reg <= i2_domand1_G4_mul0_G16_mul2_G256_inv0;
        p4_domand1_G4_mul0_G16_mul2_G256_inv0_reg <= p4_domand1_G4_mul0_G16_mul2_G256_inv0;
        z4689_assgn46890 <= z4689_assgn4689;
        z4689_assgn46891 <= z4689_assgn46890;
        z1905_assgn1905 <= z4689_assgn46891;
        z4693_assgn46930 <= z4693_assgn4693;
        z4693_assgn46931 <= z4693_assgn46930;
        z1907_assgn1907 <= z4693_assgn46931;
        z4697_assgn46970 <= z4697_assgn4697;
        z4697_assgn46971 <= z4697_assgn46970;
        z1909_assgn1909 <= z4697_assgn46971;
        z4701_assgn47010 <= z4701_assgn4701;
        z4701_assgn47011 <= z4701_assgn47010;
        z1911_assgn1911 <= z4701_assgn47011;
        z4705_assgn47050 <= z4705_assgn4705;
        z4705_assgn47051 <= z4705_assgn47050;
        z1913_assgn1913 <= z4705_assgn47051;
        z4709_assgn47090 <= z4709_assgn4709;
        z4709_assgn47091 <= z4709_assgn47090;
        z1915_assgn1915 <= z4709_assgn47091;
        i1_domand2_G4_mul0_G16_mul2_G256_inv0_reg <= i1_domand2_G4_mul0_G16_mul2_G256_inv0;
        p1_domand2_G4_mul0_G16_mul2_G256_inv0_reg <= p1_domand2_G4_mul0_G16_mul2_G256_inv0;
        i2_domand2_G4_mul0_G16_mul2_G256_inv0_reg <= i2_domand2_G4_mul0_G16_mul2_G256_inv0;
        p4_domand2_G4_mul0_G16_mul2_G256_inv0_reg <= p4_domand2_G4_mul0_G16_mul2_G256_inv0;
        z4721_assgn47210 <= z4721_assgn4721;
        z4721_assgn47211 <= z4721_assgn47210;
        z4721_assgn47212 <= z4721_assgn47211;
        z1925_assgn1925 <= z4721_assgn47212;
        z4725_assgn47250 <= z4725_assgn4725;
        z4725_assgn47251 <= z4725_assgn47250;
        z4725_assgn47252 <= z4725_assgn47251;
        z1927_assgn1927 <= z4725_assgn47252;
        z4733_assgn47330 <= z4733_assgn4733;
        z4733_assgn47331 <= z4733_assgn47330;
        z4733_assgn47332 <= z4733_assgn47331;
        z1933_assgn1933 <= z4733_assgn47332;
        z4737_assgn47370 <= z4737_assgn4737;
        z4737_assgn47371 <= z4737_assgn47370;
        z4737_assgn47372 <= z4737_assgn47371;
        z1935_assgn1935 <= z4737_assgn47372;
        z4741_assgn47410 <= z4741_assgn4741;
        z4741_assgn47411 <= z4741_assgn47410;
        z4741_assgn47412 <= z4741_assgn47411;
        z1937_assgn1937 <= z4741_assgn47412;
        z4745_assgn47450 <= z4745_assgn4745;
        z4745_assgn47451 <= z4745_assgn47450;
        z4745_assgn47452 <= z4745_assgn47451;
        z1939_assgn1939 <= z4745_assgn47452;
        z4749_assgn47490 <= z4749_assgn4749;
        z4749_assgn47491 <= z4749_assgn47490;
        z4749_assgn47492 <= z4749_assgn47491;
        z1941_assgn1941 <= z4749_assgn47492;
        z4753_assgn47530 <= z4753_assgn4753;
        z4753_assgn47531 <= z4753_assgn47530;
        z4753_assgn47532 <= z4753_assgn47531;
        z1943_assgn1943 <= z4753_assgn47532;
        z4765_assgn47650 <= z4765_assgn4765;
        z4765_assgn47651 <= z4765_assgn47650;
        z4765_assgn47652 <= z4765_assgn47651;
        z1953_assgn1953 <= z4765_assgn47652;
        z4769_assgn47690 <= z4769_assgn4769;
        z4769_assgn47691 <= z4769_assgn47690;
        z4769_assgn47692 <= z4769_assgn47691;
        z1955_assgn1955 <= z4769_assgn47692;
        z4783_assgn47830 <= z4783_assgn4783;
        z4783_assgn47831 <= z4783_assgn47830;
        z1967_assgn1967 <= z4783_assgn47831;
        z4787_assgn47870 <= z4787_assgn4787;
        z4787_assgn47871 <= z4787_assgn47870;
        z1969_assgn1969 <= z4787_assgn47871;
        z4791_assgn47910 <= z4791_assgn4791;
        z4791_assgn47911 <= z4791_assgn47910;
        z1971_assgn1971 <= z4791_assgn47911;
        z4795_assgn47950 <= z4795_assgn4795;
        z4795_assgn47951 <= z4795_assgn47950;
        z1973_assgn1973 <= z4795_assgn47951;
        z4799_assgn47990 <= z4799_assgn4799;
        z4799_assgn47991 <= z4799_assgn47990;
        z1975_assgn1975 <= z4799_assgn47991;
        z4803_assgn48030 <= z4803_assgn4803;
        z4803_assgn48031 <= z4803_assgn48030;
        z1977_assgn1977 <= z4803_assgn48031;
        z4829_assgn48290 <= z4829_assgn4829;
        z4829_assgn48291 <= z4829_assgn48290;
        z2001_assgn2001 <= z4829_assgn48291;
        z4833_assgn48330 <= z4833_assgn4833;
        z4833_assgn48331 <= z4833_assgn48330;
        z2003_assgn2003 <= z4833_assgn48331;
        z4837_assgn48370 <= z4837_assgn4837;
        z4837_assgn48371 <= z4837_assgn48370;
        z2005_assgn2005 <= z4837_assgn48371;
        z4841_assgn48410 <= z4841_assgn4841;
        z4841_assgn48411 <= z4841_assgn48410;
        z2007_assgn2007 <= z4841_assgn48411;
        z4845_assgn48450 <= z4845_assgn4845;
        z4845_assgn48451 <= z4845_assgn48450;
        z2009_assgn2009 <= z4845_assgn48451;
        z4849_assgn48490 <= z4849_assgn4849;
        z4849_assgn48491 <= z4849_assgn48490;
        z2011_assgn2011 <= z4849_assgn48491;
        i1_domand0_G4_mul1_G16_mul2_G256_inv0_reg <= i1_domand0_G4_mul1_G16_mul2_G256_inv0;
        p1_domand0_G4_mul1_G16_mul2_G256_inv0_reg <= p1_domand0_G4_mul1_G16_mul2_G256_inv0;
        i2_domand0_G4_mul1_G16_mul2_G256_inv0_reg <= i2_domand0_G4_mul1_G16_mul2_G256_inv0;
        p4_domand0_G4_mul1_G16_mul2_G256_inv0_reg <= p4_domand0_G4_mul1_G16_mul2_G256_inv0;
        z4859_assgn48590 <= z4859_assgn4859;
        z4859_assgn48591 <= z4859_assgn48590;
        z2019_assgn2019 <= z4859_assgn48591;
        z4863_assgn48630 <= z4863_assgn4863;
        z4863_assgn48631 <= z4863_assgn48630;
        z2021_assgn2021 <= z4863_assgn48631;
        z4867_assgn48670 <= z4867_assgn4867;
        z4867_assgn48671 <= z4867_assgn48670;
        z2023_assgn2023 <= z4867_assgn48671;
        z4871_assgn48710 <= z4871_assgn4871;
        z4871_assgn48711 <= z4871_assgn48710;
        z2025_assgn2025 <= z4871_assgn48711;
        z4875_assgn48750 <= z4875_assgn4875;
        z4875_assgn48751 <= z4875_assgn48750;
        z2027_assgn2027 <= z4875_assgn48751;
        z4879_assgn48790 <= z4879_assgn4879;
        z4879_assgn48791 <= z4879_assgn48790;
        z2029_assgn2029 <= z4879_assgn48791;
        i1_domand1_G4_mul1_G16_mul2_G256_inv0_reg <= i1_domand1_G4_mul1_G16_mul2_G256_inv0;
        p1_domand1_G4_mul1_G16_mul2_G256_inv0_reg <= p1_domand1_G4_mul1_G16_mul2_G256_inv0;
        i2_domand1_G4_mul1_G16_mul2_G256_inv0_reg <= i2_domand1_G4_mul1_G16_mul2_G256_inv0;
        p4_domand1_G4_mul1_G16_mul2_G256_inv0_reg <= p4_domand1_G4_mul1_G16_mul2_G256_inv0;
        z4893_assgn48930 <= z4893_assgn4893;
        z4893_assgn48931 <= z4893_assgn48930;
        z2041_assgn2041 <= z4893_assgn48931;
        z4897_assgn48970 <= z4897_assgn4897;
        z4897_assgn48971 <= z4897_assgn48970;
        z2043_assgn2043 <= z4897_assgn48971;
        z4901_assgn49010 <= z4901_assgn4901;
        z4901_assgn49011 <= z4901_assgn49010;
        z2045_assgn2045 <= z4901_assgn49011;
        z4905_assgn49050 <= z4905_assgn4905;
        z4905_assgn49051 <= z4905_assgn49050;
        z2047_assgn2047 <= z4905_assgn49051;
        z4909_assgn49090 <= z4909_assgn4909;
        z4909_assgn49091 <= z4909_assgn49090;
        z2049_assgn2049 <= z4909_assgn49091;
        z4913_assgn49130 <= z4913_assgn4913;
        z4913_assgn49131 <= z4913_assgn49130;
        z2051_assgn2051 <= z4913_assgn49131;
        i1_domand2_G4_mul1_G16_mul2_G256_inv0_reg <= i1_domand2_G4_mul1_G16_mul2_G256_inv0;
        p1_domand2_G4_mul1_G16_mul2_G256_inv0_reg <= p1_domand2_G4_mul1_G16_mul2_G256_inv0;
        i2_domand2_G4_mul1_G16_mul2_G256_inv0_reg <= i2_domand2_G4_mul1_G16_mul2_G256_inv0;
        p4_domand2_G4_mul1_G16_mul2_G256_inv0_reg <= p4_domand2_G4_mul1_G16_mul2_G256_inv0;
        z4925_assgn49250 <= z4925_assgn4925;
        z4925_assgn49251 <= z4925_assgn49250;
        z4925_assgn49252 <= z4925_assgn49251;
        z2061_assgn2061 <= z4925_assgn49252;
        z4929_assgn49290 <= z4929_assgn4929;
        z4929_assgn49291 <= z4929_assgn49290;
        z4929_assgn49292 <= z4929_assgn49291;
        z2063_assgn2063 <= z4929_assgn49292;
        z4947_assgn49470 <= z4947_assgn4947;
        z4947_assgn49471 <= z4947_assgn49470;
        z2079_assgn2079 <= z4947_assgn49471;
        z4951_assgn49510 <= z4951_assgn4951;
        z4951_assgn49511 <= z4951_assgn49510;
        z2081_assgn2081 <= z4951_assgn49511;
        z4955_assgn49550 <= z4955_assgn4955;
        z4955_assgn49551 <= z4955_assgn49550;
        z2083_assgn2083 <= z4955_assgn49551;
        z4959_assgn49590 <= z4959_assgn4959;
        z4959_assgn49591 <= z4959_assgn49590;
        z2085_assgn2085 <= z4959_assgn49591;
        z4963_assgn49630 <= z4963_assgn4963;
        z4963_assgn49631 <= z4963_assgn49630;
        z2087_assgn2087 <= z4963_assgn49631;
        z4967_assgn49670 <= z4967_assgn4967;
        z4967_assgn49671 <= z4967_assgn49670;
        z2089_assgn2089 <= z4967_assgn49671;
        z4993_assgn49930 <= z4993_assgn4993;
        z4993_assgn49931 <= z4993_assgn49930;
        z2113_assgn2113 <= z4993_assgn49931;
        z4997_assgn49970 <= z4997_assgn4997;
        z4997_assgn49971 <= z4997_assgn49970;
        z2115_assgn2115 <= z4997_assgn49971;
        z5001_assgn50010 <= z5001_assgn5001;
        z5001_assgn50011 <= z5001_assgn50010;
        z2117_assgn2117 <= z5001_assgn50011;
        z5005_assgn50050 <= z5005_assgn5005;
        z5005_assgn50051 <= z5005_assgn50050;
        z2119_assgn2119 <= z5005_assgn50051;
        z5009_assgn50090 <= z5009_assgn5009;
        z5009_assgn50091 <= z5009_assgn50090;
        z2121_assgn2121 <= z5009_assgn50091;
        z5013_assgn50130 <= z5013_assgn5013;
        z5013_assgn50131 <= z5013_assgn50130;
        z2123_assgn2123 <= z5013_assgn50131;
        i1_domand0_G4_mul2_G16_mul2_G256_inv0_reg <= i1_domand0_G4_mul2_G16_mul2_G256_inv0;
        p1_domand0_G4_mul2_G16_mul2_G256_inv0_reg <= p1_domand0_G4_mul2_G16_mul2_G256_inv0;
        i2_domand0_G4_mul2_G16_mul2_G256_inv0_reg <= i2_domand0_G4_mul2_G16_mul2_G256_inv0;
        p4_domand0_G4_mul2_G16_mul2_G256_inv0_reg <= p4_domand0_G4_mul2_G16_mul2_G256_inv0;
        z5023_assgn50230 <= z5023_assgn5023;
        z5023_assgn50231 <= z5023_assgn50230;
        z2131_assgn2131 <= z5023_assgn50231;
        z5027_assgn50270 <= z5027_assgn5027;
        z5027_assgn50271 <= z5027_assgn50270;
        z2133_assgn2133 <= z5027_assgn50271;
        z5031_assgn50310 <= z5031_assgn5031;
        z5031_assgn50311 <= z5031_assgn50310;
        z2135_assgn2135 <= z5031_assgn50311;
        z5035_assgn50350 <= z5035_assgn5035;
        z5035_assgn50351 <= z5035_assgn50350;
        z2137_assgn2137 <= z5035_assgn50351;
        z5039_assgn50390 <= z5039_assgn5039;
        z5039_assgn50391 <= z5039_assgn50390;
        z2139_assgn2139 <= z5039_assgn50391;
        z5043_assgn50430 <= z5043_assgn5043;
        z5043_assgn50431 <= z5043_assgn50430;
        z2141_assgn2141 <= z5043_assgn50431;
        i1_domand1_G4_mul2_G16_mul2_G256_inv0_reg <= i1_domand1_G4_mul2_G16_mul2_G256_inv0;
        p1_domand1_G4_mul2_G16_mul2_G256_inv0_reg <= p1_domand1_G4_mul2_G16_mul2_G256_inv0;
        i2_domand1_G4_mul2_G16_mul2_G256_inv0_reg <= i2_domand1_G4_mul2_G16_mul2_G256_inv0;
        p4_domand1_G4_mul2_G16_mul2_G256_inv0_reg <= p4_domand1_G4_mul2_G16_mul2_G256_inv0;
        z5057_assgn50570 <= z5057_assgn5057;
        z5057_assgn50571 <= z5057_assgn50570;
        z2153_assgn2153 <= z5057_assgn50571;
        z5061_assgn50610 <= z5061_assgn5061;
        z5061_assgn50611 <= z5061_assgn50610;
        z2155_assgn2155 <= z5061_assgn50611;
        z5065_assgn50650 <= z5065_assgn5065;
        z5065_assgn50651 <= z5065_assgn50650;
        z2157_assgn2157 <= z5065_assgn50651;
        z5069_assgn50690 <= z5069_assgn5069;
        z5069_assgn50691 <= z5069_assgn50690;
        z2159_assgn2159 <= z5069_assgn50691;
        z5073_assgn50730 <= z5073_assgn5073;
        z5073_assgn50731 <= z5073_assgn50730;
        z2161_assgn2161 <= z5073_assgn50731;
        z5077_assgn50770 <= z5077_assgn5077;
        z5077_assgn50771 <= z5077_assgn50770;
        z2163_assgn2163 <= z5077_assgn50771;
        i1_domand2_G4_mul2_G16_mul2_G256_inv0_reg <= i1_domand2_G4_mul2_G16_mul2_G256_inv0;
        p1_domand2_G4_mul2_G16_mul2_G256_inv0_reg <= p1_domand2_G4_mul2_G16_mul2_G256_inv0;
        i2_domand2_G4_mul2_G16_mul2_G256_inv0_reg <= i2_domand2_G4_mul2_G16_mul2_G256_inv0;
        p4_domand2_G4_mul2_G16_mul2_G256_inv0_reg <= p4_domand2_G4_mul2_G16_mul2_G256_inv0;
        z5089_assgn50890 <= z5089_assgn5089;
        z5089_assgn50891 <= z5089_assgn50890;
        z5089_assgn50892 <= z5089_assgn50891;
        z2173_assgn2173 <= z5089_assgn50892;
        z5093_assgn50930 <= z5093_assgn5093;
        z5093_assgn50931 <= z5093_assgn50930;
        z5093_assgn50932 <= z5093_assgn50931;
        z2175_assgn2175 <= z5093_assgn50932;
        z5105_assgn51050 <= z5105_assgn5105;
        z5105_assgn51051 <= z5105_assgn51050;
        z5105_assgn51052 <= z5105_assgn51051;
        z2185_assgn2185 <= z5105_assgn51052;
        z5109_assgn51090 <= z5109_assgn5109;
        z5109_assgn51091 <= z5109_assgn51090;
        z5109_assgn51092 <= z5109_assgn51091;
        z2187_assgn2187 <= z5109_assgn51092;
        z5117_assgn51170 <= z5117_assgn5117;
        z5117_assgn51171 <= z5117_assgn51170;
        z5117_assgn51172 <= z5117_assgn51171;
        z2193_assgn2193 <= z5117_assgn51172;
        z5121_assgn51210 <= z5121_assgn5121;
        z5121_assgn51211 <= z5121_assgn51210;
        z5121_assgn51212 <= z5121_assgn51211;
        z2195_assgn2195 <= z5121_assgn51212;
        z5133_assgn51330 <= z5133_assgn5133;
        z5133_assgn51331 <= z5133_assgn51330;
        z5133_assgn51332 <= z5133_assgn51331;
        z2205_assgn2205 <= z5133_assgn51332;
        z5141_assgn51410 <= z5141_assgn5141;
        z5141_assgn51411 <= z5141_assgn51410;
        z5141_assgn51412 <= z5141_assgn51411;
        z2211_assgn2211 <= z5141_assgn51412;
        z5145_assgn51450 <= z5145_assgn5145;
        z5145_assgn51451 <= z5145_assgn51450;
        z5145_assgn51452 <= z5145_assgn51451;
        z2214_assgn2214 <= z5145_assgn51452;
        z5151_assgn51510 <= z5151_assgn5151;
        z5151_assgn51511 <= z5151_assgn51510;
        z5151_assgn51512 <= z5151_assgn51511;
        z2217_assgn2217 <= z5151_assgn51512;
        z5157_assgn51570 <= z5157_assgn5157;
        z5157_assgn51571 <= z5157_assgn51570;
        z5157_assgn51572 <= z5157_assgn51571;
        z2221_assgn2221 <= z5157_assgn51572;
        z5163_assgn51630 <= z5163_assgn5163;
        z5163_assgn51631 <= z5163_assgn51630;
        z5163_assgn51632 <= z5163_assgn51631;
        z2225_assgn2225 <= z5163_assgn51632;
        z5173_assgn51730 <= z5173_assgn5173;
        z5173_assgn51731 <= z5173_assgn51730;
        z5173_assgn51732 <= z5173_assgn51731;
        z2233_assgn2233 <= z5173_assgn51732;
        z5179_assgn51790 <= z5179_assgn5179;
        z5179_assgn51791 <= z5179_assgn51790;
        z5179_assgn51792 <= z5179_assgn51791;
        z2237_assgn2237 <= z5179_assgn51792;
        z5185_assgn51850 <= z5185_assgn5185;
        z5185_assgn51851 <= z5185_assgn51850;
        z5185_assgn51852 <= z5185_assgn51851;
        z2241_assgn2241 <= z5185_assgn51852;
        z5195_assgn51950 <= z5195_assgn5195;
        z5195_assgn51951 <= z5195_assgn51950;
        z5195_assgn51952 <= z5195_assgn51951;
        z2249_assgn2249 <= z5195_assgn51952;
        z5201_assgn52010 <= z5201_assgn5201;
        z5201_assgn52011 <= z5201_assgn52010;
        z5201_assgn52012 <= z5201_assgn52011;
        z2253_assgn2253 <= z5201_assgn52012;
        z5207_assgn52070 <= z5207_assgn5207;
        z5207_assgn52071 <= z5207_assgn52070;
        z5207_assgn52072 <= z5207_assgn52071;
        z2257_assgn2257 <= z5207_assgn52072;
        z5217_assgn52170 <= z5217_assgn5217;
        z5217_assgn52171 <= z5217_assgn52170;
        z5217_assgn52172 <= z5217_assgn52171;
        z2265_assgn2265 <= z5217_assgn52172;
        z5223_assgn52230 <= z5223_assgn5223;
        z5223_assgn52231 <= z5223_assgn52230;
        z5223_assgn52232 <= z5223_assgn52231;
        z2269_assgn2269 <= z5223_assgn52232;
        z5229_assgn52290 <= z5229_assgn5229;
        z5229_assgn52291 <= z5229_assgn52290;
        z5229_assgn52292 <= z5229_assgn52291;
        z2273_assgn2273 <= z5229_assgn52292;
        z5239_assgn52390 <= z5239_assgn5239;
        z5239_assgn52391 <= z5239_assgn52390;
        z5239_assgn52392 <= z5239_assgn52391;
        z2281_assgn2281 <= z5239_assgn52392;
        z5245_assgn52450 <= z5245_assgn5245;
        z5245_assgn52451 <= z5245_assgn52450;
        z5245_assgn52452 <= z5245_assgn52451;
        z2285_assgn2285 <= z5245_assgn52452;
        z5251_assgn52510 <= z5251_assgn5251;
        z5251_assgn52511 <= z5251_assgn52510;
        z5251_assgn52512 <= z5251_assgn52511;
        z2289_assgn2289 <= z5251_assgn52512;
        z5261_assgn52610 <= z5261_assgn5261;
        z5261_assgn52611 <= z5261_assgn52610;
        z5261_assgn52612 <= z5261_assgn52611;
        z2297_assgn2297 <= z5261_assgn52612;
        z5267_assgn52670 <= z5267_assgn5267;
        z5267_assgn52671 <= z5267_assgn52670;
        z5267_assgn52672 <= z5267_assgn52671;
        z2301_assgn2301 <= z5267_assgn52672;
        z5273_assgn52730 <= z5273_assgn5273;
        z5273_assgn52731 <= z5273_assgn52730;
        z5273_assgn52732 <= z5273_assgn52731;
        z2305_assgn2305 <= z5273_assgn52732;
        z5283_assgn52830 <= z5283_assgn5283;
        z5283_assgn52831 <= z5283_assgn52830;
        z5283_assgn52832 <= z5283_assgn52831;
        z2313_assgn2313 <= z5283_assgn52832;
        z5289_assgn52890 <= z5289_assgn5289;
        z5289_assgn52891 <= z5289_assgn52890;
        z5289_assgn52892 <= z5289_assgn52891;
        z2317_assgn2317 <= z5289_assgn52892;
        z5295_assgn52950 <= z5295_assgn5295;
        z5295_assgn52951 <= z5295_assgn52950;
        z5295_assgn52952 <= z5295_assgn52951;
        z2321_assgn2321 <= z5295_assgn52952;
        z5305_assgn53050 <= z5305_assgn5305;
        z5305_assgn53051 <= z5305_assgn53050;
        z5305_assgn53052 <= z5305_assgn53051;
        z2329_assgn2329 <= z5305_assgn53052;
        z5315_assgn53150 <= z5315_assgn5315;
        z5315_assgn53151 <= z5315_assgn53150;
        z5315_assgn53152 <= z5315_assgn53151;
        z2337_assgn2337 <= z5315_assgn53152;
        z5323_assgn53230 <= z5323_assgn5323;
        z5323_assgn53231 <= z5323_assgn53230;
        z5323_assgn53232 <= z5323_assgn53231;
        z2343_assgn2343 <= z5323_assgn53232;
        z5327_assgn53270 <= z5327_assgn5327;
        z5327_assgn53271 <= z5327_assgn53270;
        z5327_assgn53272 <= z5327_assgn53271;
        z2346_assgn2346 <= z5327_assgn53272;
        z5333_assgn53330 <= z5333_assgn5333;
        z5333_assgn53331 <= z5333_assgn53330;
        z5333_assgn53332 <= z5333_assgn53331;
        z2349_assgn2349 <= z5333_assgn53332;
        z5339_assgn53390 <= z5339_assgn5339;
        z5339_assgn53391 <= z5339_assgn53390;
        z5339_assgn53392 <= z5339_assgn53391;
        z2353_assgn2353 <= z5339_assgn53392;
        z5345_assgn53450 <= z5345_assgn5345;
        z5345_assgn53451 <= z5345_assgn53450;
        z5345_assgn53452 <= z5345_assgn53451;
        z2357_assgn2357 <= z5345_assgn53452;
        z5355_assgn53550 <= z5355_assgn5355;
        z5355_assgn53551 <= z5355_assgn53550;
        z5355_assgn53552 <= z5355_assgn53551;
        z2365_assgn2365 <= z5355_assgn53552;
        z5361_assgn53610 <= z5361_assgn5361;
        z5361_assgn53611 <= z5361_assgn53610;
        z5361_assgn53612 <= z5361_assgn53611;
        z2369_assgn2369 <= z5361_assgn53612;
        z5367_assgn53670 <= z5367_assgn5367;
        z5367_assgn53671 <= z5367_assgn53670;
        z5367_assgn53672 <= z5367_assgn53671;
        z2373_assgn2373 <= z5367_assgn53672;
        z5377_assgn53770 <= z5377_assgn5377;
        z5377_assgn53771 <= z5377_assgn53770;
        z5377_assgn53772 <= z5377_assgn53771;
        z2381_assgn2381 <= z5377_assgn53772;
        z5383_assgn53830 <= z5383_assgn5383;
        z5383_assgn53831 <= z5383_assgn53830;
        z5383_assgn53832 <= z5383_assgn53831;
        z2385_assgn2385 <= z5383_assgn53832;
        z5389_assgn53890 <= z5389_assgn5389;
        z5389_assgn53891 <= z5389_assgn53890;
        z5389_assgn53892 <= z5389_assgn53891;
        z2389_assgn2389 <= z5389_assgn53892;
        z5399_assgn53990 <= z5399_assgn5399;
        z5399_assgn53991 <= z5399_assgn53990;
        z5399_assgn53992 <= z5399_assgn53991;
        z2397_assgn2397 <= z5399_assgn53992;
        z5405_assgn54050 <= z5405_assgn5405;
        z5405_assgn54051 <= z5405_assgn54050;
        z5405_assgn54052 <= z5405_assgn54051;
        z2401_assgn2401 <= z5405_assgn54052;
        z5411_assgn54110 <= z5411_assgn5411;
        z5411_assgn54111 <= z5411_assgn54110;
        z5411_assgn54112 <= z5411_assgn54111;
        z2405_assgn2405 <= z5411_assgn54112;
        z5421_assgn54210 <= z5421_assgn5421;
        z5421_assgn54211 <= z5421_assgn54210;
        z5421_assgn54212 <= z5421_assgn54211;
        z2413_assgn2413 <= z5421_assgn54212;
        z5427_assgn54270 <= z5427_assgn5427;
        z5427_assgn54271 <= z5427_assgn54270;
        z5427_assgn54272 <= z5427_assgn54271;
        z2417_assgn2417 <= z5427_assgn54272;
        z5433_assgn54330 <= z5433_assgn5433;
        z5433_assgn54331 <= z5433_assgn54330;
        z5433_assgn54332 <= z5433_assgn54331;
        z2421_assgn2421 <= z5433_assgn54332;
        z5443_assgn54430 <= z5443_assgn5443;
        z5443_assgn54431 <= z5443_assgn54430;
        z5443_assgn54432 <= z5443_assgn54431;
        z2429_assgn2429 <= z5443_assgn54432;
        z5449_assgn54490 <= z5449_assgn5449;
        z5449_assgn54491 <= z5449_assgn54490;
        z5449_assgn54492 <= z5449_assgn54491;
        z2433_assgn2433 <= z5449_assgn54492;
        z5455_assgn54550 <= z5455_assgn5455;
        z5455_assgn54551 <= z5455_assgn54550;
        z5455_assgn54552 <= z5455_assgn54551;
        z2437_assgn2437 <= z5455_assgn54552;
        z5465_assgn54650 <= z5465_assgn5465;
        z5465_assgn54651 <= z5465_assgn54650;
        z5465_assgn54652 <= z5465_assgn54651;
        z2445_assgn2445 <= z5465_assgn54652;
        z5471_assgn54710 <= z5471_assgn5471;
        z5471_assgn54711 <= z5471_assgn54710;
        z5471_assgn54712 <= z5471_assgn54711;
        z2449_assgn2449 <= z5471_assgn54712;
        z5477_assgn54770 <= z5477_assgn5477;
        z5477_assgn54771 <= z5477_assgn54770;
        z5477_assgn54772 <= z5477_assgn54771;
        z2453_assgn2453 <= z5477_assgn54772;
        z5487_assgn54870 <= z5487_assgn5487;
        z5487_assgn54871 <= z5487_assgn54870;
        z5487_assgn54872 <= z5487_assgn54871;
        z2461_assgn2461 <= z5487_assgn54872;
        z5493_assgn54930 <= z5493_assgn5493;
        z5493_assgn54931 <= z5493_assgn54930;
        z5493_assgn54932 <= z5493_assgn54931;
        z2465_assgn2465 <= z5493_assgn54932;
        y0 <= (t6 ^ z2465_assgn2465);
        y1 <= t7;
    end

endmodule



        