module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    reg z5_assgn5;
    wire z275_assgn275;
    reg z275_assgn2750;
    reg x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    reg z7_assgn7;
    wire z285_assgn285;
    reg z285_assgn2850;
    reg x3_1_inp;
    wire r_inp;
    reg x1_0_inp_reg;
    wire L0_0;
    wire L1_0;
    wire z293_assgn293;
    reg z293_assgn2930;
    reg z293_assgn2931;
    reg z293_assgn2932;
    reg z47_assgn47;
    wire z295_assgn295;
    reg z295_assgn2950;
    reg z295_assgn2951;
    reg z48_assgn48;
    wire L8_0;
    wire z299_assgn299;
    reg z299_assgn2990;
    reg z50_assgn50;
    wire L5_0;
    reg x1_1_inp_reg;
    wire L0_1;
    wire L1_1;
    wire z307_assgn307;
    reg z307_assgn3070;
    reg z307_assgn3071;
    reg z307_assgn3072;
    reg z55_assgn55;
    wire z309_assgn309;
    reg z309_assgn3090;
    reg z309_assgn3091;
    reg z56_assgn56;
    wire L8_1;
    wire z313_assgn313;
    reg z313_assgn3130;
    reg z58_assgn58;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire z333_assgn333;
    reg z333_assgn3330;
    reg z75_assgn75;
    wire z335_assgn335;
    reg z335_assgn3350;
    reg z335_assgn3351;
    reg z76_assgn76;
    wire L2_0;
    wire z339_assgn339;
    reg z339_assgn3390;
    reg z78_assgn78;
    reg x3_0_inp_reg;
    wire L3_0;
    wire z343_assgn343;
    reg z343_assgn3430;
    reg z79_assgn79;
    wire z345_assgn345;
    reg z345_assgn3450;
    reg z345_assgn3451;
    reg z80_assgn80;
    wire L2_1;
    wire z349_assgn349;
    reg z349_assgn3490;
    reg z82_assgn82;
    reg x3_1_inp_reg;
    wire L3_1;
    wire a0_neg_hpc20;
    wire a1_neg_hpc20;
    reg r_inp_reg;
    wire u0_hpc20;
    wire u1_hpc20;
    wire v0_hpc20;
    wire v1_hpc20;
    reg Q1_0_reg;
    wire p0_hpc20;
    reg v1_hpc20_reg;
    wire p1_hpc20;
    reg u0_hpc20_reg;
    reg p1_hpc20_reg;
    wire p01_hpc20;
    reg p0_hpc20_reg;
    wire T0_0;
    reg Q1_1_reg;
    wire p2_hpc20;
    reg v0_hpc20_reg;
    wire p3_hpc20;
    reg u1_hpc20_reg;
    reg p3_hpc20_reg;
    wire p23_hpc20;
    reg p2_hpc20_reg;
    wire T0_1;
    wire z1_assgn1;
    reg L10_0;
    wire z2_assgn2;
    reg L10_1;
    wire z3_assgn3;
    wire z391_assgn391;
    reg z391_assgn3910;
    reg a0_neg_hpc21;
    wire z4_assgn4;
    wire z395_assgn395;
    reg z395_assgn3950;
    reg a1_neg_hpc21;
    wire z397_assgn397;
    reg z397_assgn3970;
    reg z127_assgn127;
    wire u0_hpc21;
    wire z401_assgn401;
    reg z401_assgn4010;
    reg z129_assgn129;
    wire u1_hpc21;
    wire v0_hpc21;
    wire v1_hpc21;
    wire z409_assgn409;
    reg z409_assgn4090;
    reg z136_assgn136;
    reg Q4_0_reg;
    wire p0_hpc21;
    wire z413_assgn413;
    reg z413_assgn4130;
    reg z138_assgn138;
    reg v1_hpc21_reg;
    wire p1_hpc21;
    reg u0_hpc21_reg;
    reg p1_hpc21_reg;
    wire p01_hpc21;
    reg p0_hpc21_reg;
    wire T2_0;
    wire z421_assgn421;
    reg z421_assgn4210;
    reg z144_assgn144;
    reg Q4_1_reg;
    wire p2_hpc21;
    wire z425_assgn425;
    reg z425_assgn4250;
    reg z146_assgn146;
    reg v0_hpc21_reg;
    wire p3_hpc21;
    reg u1_hpc21_reg;
    reg p3_hpc21_reg;
    wire p23_hpc21;
    reg p2_hpc21_reg;
    wire T2_1;
    reg T0_0_reg;
    wire Q2_0;
    wire L4_0;
    wire Q7_0;
    wire Q6_0;
    reg T0_1_reg;
    wire Q2_1;
    wire L4_1;
    wire Q7_1;
    wire Q6_1;
    wire a0_neg_hpc22;
    wire a1_neg_hpc22;
    wire z453_assgn453;
    reg z453_assgn4530;
    reg z453_assgn4531;
    reg z171_assgn171;
    wire u0_hpc22;
    wire z457_assgn457;
    reg z457_assgn4570;
    reg z457_assgn4571;
    reg z173_assgn173;
    wire u1_hpc22;
    wire z461_assgn461;
    reg z461_assgn4610;
    reg z175_assgn175;
    wire v0_hpc22;
    wire z465_assgn465;
    reg z465_assgn4650;
    reg z177_assgn177;
    wire v1_hpc22;
    reg Q3_0_reg;
    wire p0_hpc22;
    reg v1_hpc22_reg;
    wire p1_hpc22;
    reg u0_hpc22_reg;
    reg p1_hpc22_reg;
    wire p01_hpc22;
    reg p0_hpc22_reg;
    wire T1_0;
    reg Q3_1_reg;
    wire p2_hpc22;
    reg v0_hpc22_reg;
    wire p3_hpc22;
    reg u1_hpc22_reg;
    reg p3_hpc22_reg;
    wire p23_hpc22;
    reg p2_hpc22_reg;
    wire T1_1;
    wire a0_neg_hpc23;
    wire a1_neg_hpc23;
    wire z489_assgn489;
    reg z489_assgn4890;
    reg z489_assgn4891;
    reg z199_assgn199;
    wire u0_hpc23;
    wire z493_assgn493;
    reg z493_assgn4930;
    reg z493_assgn4931;
    reg z201_assgn201;
    wire u1_hpc23;
    wire z497_assgn497;
    reg z497_assgn4970;
    reg z203_assgn203;
    wire v0_hpc23;
    wire z501_assgn501;
    reg z501_assgn5010;
    reg z205_assgn205;
    wire v1_hpc23;
    reg Q7_0_reg;
    wire p0_hpc23;
    reg v1_hpc23_reg;
    wire p1_hpc23;
    reg u0_hpc23_reg;
    reg p1_hpc23_reg;
    wire p01_hpc23;
    reg p0_hpc23_reg;
    wire T3_0;
    reg Q7_1_reg;
    wire p2_hpc23;
    reg v0_hpc23_reg;
    wire p3_hpc23;
    reg u1_hpc23_reg;
    reg p3_hpc23_reg;
    wire p23_hpc23;
    reg p2_hpc23_reg;
    wire T3_1;
    wire z521_assgn521;
    reg z521_assgn5210;
    reg z224_assgn224;
    wire L7_0;
    wire L11_0;
    wire z527_assgn527;
    reg z527_assgn5270;
    reg z228_assgn228;
    wire L7_1;
    wire L11_1;
    reg T2_0_reg;
    wire Y0_01;
    wire Y1_01;
    reg T2_1_reg;
    wire Y0_11;
    wire Y1_11;
    wire z541_assgn541;
    reg z541_assgn5410;
    reg z240_assgn240;
    wire z9_assgn9;
    wire z11_assgn11;
    wire z553_assgn553;
    reg z553_assgn5530;
    reg z249_assgn249;
    wire z13_assgn13;
    wire z559_assgn559;
    reg z559_assgn5590;
    reg z254_assgn254;
    wire z15_assgn15;
    wire z17_assgn17;
    wire z571_assgn571;
    reg z571_assgn5710;
    reg z263_assgn263;
    wire z19_assgn19;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign z275_assgn275 = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign z285_assgn285 = x3_1;
    assign r_inp = r;
    assign L0_0 = (x1_0_inp_reg ^ z5_assgn5);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign z293_assgn293 = x0_0_inp;
    assign z295_assgn295 = z5_assgn5;
    assign L8_0 = (z48_assgn48 ^ z47_assgn47);
    assign z299_assgn299 = x0_0_inp;
    assign L5_0 = (z50_assgn50 ^ x3_0_inp);
    assign L0_1 = (x1_1_inp_reg ^ z7_assgn7);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign z307_assgn307 = x0_1_inp;
    assign z309_assgn309 = z7_assgn7;
    assign L8_1 = (z56_assgn56 ^ z55_assgn55);
    assign z313_assgn313 = x0_1_inp;
    assign L5_1 = (z58_assgn58 ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !z5_assgn5;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !z7_assgn7;
    assign z333_assgn333 = z5_assgn5;
    assign z335_assgn335 = Q1_0;
    assign L2_0 = (z76_assgn76 ^ z75_assgn75);
    assign z339_assgn339 = Q0_0;
    assign L3_0 = (z78_assgn78 ^ x3_0_inp_reg);
    assign z343_assgn343 = z7_assgn7;
    assign z345_assgn345 = Q1_1;
    assign L2_1 = (z80_assgn80 ^ z79_assgn79);
    assign z349_assgn349 = Q0_1;
    assign L3_1 = (z82_assgn82 ^ x3_1_inp_reg);
    assign a0_neg_hpc20 = !Q0_0;
    assign a1_neg_hpc20 = !Q0_1;
    assign u0_hpc20 = (a0_neg_hpc20 & r_inp_reg);
    assign u1_hpc20 = (a1_neg_hpc20 & r_inp_reg);
    assign v0_hpc20 = (Q1_0 ^ r_inp);
    assign v1_hpc20 = (Q1_1 ^ r_inp);
    assign p0_hpc20 = (Q0_0 & Q1_0_reg);
    assign p1_hpc20 = (Q0_0 & v1_hpc20_reg);
    assign p01_hpc20 = (u0_hpc20_reg ^ p1_hpc20_reg);
    assign T0_0 = (p0_hpc20_reg ^ p01_hpc20);
    assign p2_hpc20 = (Q0_1 & Q1_1_reg);
    assign p3_hpc20 = (Q0_1 & v0_hpc20_reg);
    assign p23_hpc20 = (u1_hpc20_reg ^ p3_hpc20_reg);
    assign T0_1 = (p2_hpc20_reg ^ p23_hpc20);
    assign z1_assgn1 = !L2_0;
    assign z2_assgn2 = !L2_1;
    assign z3_assgn3 = !x1_0_inp;
    assign z391_assgn391 = z3_assgn3;
    assign z4_assgn4 = !x1_1_inp;
    assign z395_assgn395 = z4_assgn4;
    assign z397_assgn397 = r_inp;
    assign u0_hpc21 = (a0_neg_hpc21 & z127_assgn127);
    assign z401_assgn401 = r_inp;
    assign u1_hpc21 = (a1_neg_hpc21 & z129_assgn129);
    assign v0_hpc21 = (Q4_0 ^ r_inp_reg);
    assign v1_hpc21 = (Q4_1 ^ r_inp_reg);
    assign z409_assgn409 = x1_0_inp;
    assign p0_hpc21 = (z136_assgn136 & Q4_0_reg);
    assign z413_assgn413 = x1_0_inp;
    assign p1_hpc21 = (z138_assgn138 & v1_hpc21_reg);
    assign p01_hpc21 = (u0_hpc21_reg ^ p1_hpc21_reg);
    assign T2_0 = (p0_hpc21_reg ^ p01_hpc21);
    assign z421_assgn421 = x1_1_inp;
    assign p2_hpc21 = (z144_assgn144 & Q4_1_reg);
    assign z425_assgn425 = x1_1_inp;
    assign p3_hpc21 = (z146_assgn146 & v0_hpc21_reg);
    assign p23_hpc21 = (u1_hpc21_reg ^ p3_hpc21_reg);
    assign T2_1 = (p2_hpc21_reg ^ p23_hpc21);
    assign Q2_0 = (T0_0_reg ^ L2_0);
    assign L4_0 = (T0_0_reg ^ T2_0);
    assign Q7_0 = (T0_0 ^ L5_0);
    assign Q6_0 = (L4_0 ^ L3_0);
    assign Q2_1 = (T0_1_reg ^ L2_1);
    assign L4_1 = (T0_1_reg ^ T2_1);
    assign Q7_1 = (T0_1 ^ L5_1);
    assign Q6_1 = (L4_1 ^ L3_1);
    assign a0_neg_hpc22 = !Q2_0;
    assign a1_neg_hpc22 = !Q2_1;
    assign z453_assgn453 = r_inp;
    assign u0_hpc22 = (a0_neg_hpc22 & z171_assgn171);
    assign z457_assgn457 = r_inp;
    assign u1_hpc22 = (a1_neg_hpc22 & z173_assgn173);
    assign z461_assgn461 = r_inp;
    assign v0_hpc22 = (Q3_0 ^ z175_assgn175);
    assign z465_assgn465 = r_inp;
    assign v1_hpc22 = (Q3_1 ^ z177_assgn177);
    assign p0_hpc22 = (Q2_0 & Q3_0_reg);
    assign p1_hpc22 = (Q2_0 & v1_hpc22_reg);
    assign p01_hpc22 = (u0_hpc22_reg ^ p1_hpc22_reg);
    assign T1_0 = (p0_hpc22_reg ^ p01_hpc22);
    assign p2_hpc22 = (Q2_1 & Q3_1_reg);
    assign p3_hpc22 = (Q2_1 & v0_hpc22_reg);
    assign p23_hpc22 = (u1_hpc22_reg ^ p3_hpc22_reg);
    assign T1_1 = (p2_hpc22_reg ^ p23_hpc22);
    assign a0_neg_hpc23 = !Q6_0;
    assign a1_neg_hpc23 = !Q6_1;
    assign z489_assgn489 = r_inp;
    assign u0_hpc23 = (a0_neg_hpc23 & z199_assgn199);
    assign z493_assgn493 = r_inp;
    assign u1_hpc23 = (a1_neg_hpc23 & z201_assgn201);
    assign z497_assgn497 = r_inp;
    assign v0_hpc23 = (Q7_0 ^ z203_assgn203);
    assign z501_assgn501 = r_inp;
    assign v1_hpc23 = (Q7_1 ^ z205_assgn205);
    assign p0_hpc23 = (Q6_0 & Q7_0_reg);
    assign p1_hpc23 = (Q6_0 & v1_hpc23_reg);
    assign p01_hpc23 = (u0_hpc23_reg ^ p1_hpc23_reg);
    assign T3_0 = (p0_hpc23_reg ^ p01_hpc23);
    assign p2_hpc23 = (Q6_1 & Q7_1_reg);
    assign p3_hpc23 = (Q6_1 & v0_hpc23_reg);
    assign p23_hpc23 = (u1_hpc23_reg ^ p3_hpc23_reg);
    assign T3_1 = (p2_hpc23_reg ^ p23_hpc23);
    assign z521_assgn521 = T0_0;
    assign L7_0 = (z224_assgn224 ^ T1_0);
    assign L11_0 = (T1_0 ^ L10_0);
    assign z527_assgn527 = T0_1;
    assign L7_1 = (z228_assgn228 ^ T1_1);
    assign L11_1 = (T1_1 ^ L10_1);
    assign Y0_01 = (L7_0 ^ T2_0_reg);
    assign Y1_01 = (L8_0 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1_reg);
    assign Y1_11 = (L8_1 ^ T3_1);
    assign z541_assgn541 = x3_0_inp;
    assign z9_assgn9 = (z240_assgn240 ^ Y0_01);
    assign z11_assgn11 = (L11_0 ^ T2_0_reg);
    assign z553_assgn553 = L5_0;
    assign z13_assgn13 = (T2_0_reg ^ z249_assgn249);
    assign z559_assgn559 = x3_1_inp;
    assign z15_assgn15 = (z254_assgn254 ^ Y0_11);
    assign z17_assgn17 = (L11_1 ^ T2_1_reg);
    assign z571_assgn571 = L5_1;
    assign z19_assgn19 = (T2_1_reg ^ z263_assgn263);

    always @(posedge clk) begin
        z5_assgn5 <= x2_0_inp;
        z275_assgn2750 <= z275_assgn275;
        x3_0_inp <= z275_assgn2750;
        z7_assgn7 <= x2_1_inp;
        z285_assgn2850 <= z285_assgn285;
        x3_1_inp <= z285_assgn2850;
        x1_0_inp_reg <= x1_0_inp;
        z293_assgn2930 <= z293_assgn293;
        z293_assgn2931 <= z293_assgn2930;
        z293_assgn2932 <= z293_assgn2931;
        z47_assgn47 <= z293_assgn2932;
        z295_assgn2950 <= z295_assgn295;
        z295_assgn2951 <= z295_assgn2950;
        z48_assgn48 <= z295_assgn2951;
        z299_assgn2990 <= z299_assgn299;
        z50_assgn50 <= z299_assgn2990;
        x1_1_inp_reg <= x1_1_inp;
        z307_assgn3070 <= z307_assgn307;
        z307_assgn3071 <= z307_assgn3070;
        z307_assgn3072 <= z307_assgn3071;
        z55_assgn55 <= z307_assgn3072;
        z309_assgn3090 <= z309_assgn309;
        z309_assgn3091 <= z309_assgn3090;
        z56_assgn56 <= z309_assgn3091;
        z313_assgn3130 <= z313_assgn313;
        z58_assgn58 <= z313_assgn3130;
        z333_assgn3330 <= z333_assgn333;
        z75_assgn75 <= z333_assgn3330;
        z335_assgn3350 <= z335_assgn335;
        z335_assgn3351 <= z335_assgn3350;
        z76_assgn76 <= z335_assgn3351;
        z339_assgn3390 <= z339_assgn339;
        z78_assgn78 <= z339_assgn3390;
        x3_0_inp_reg <= x3_0_inp;
        z343_assgn3430 <= z343_assgn343;
        z79_assgn79 <= z343_assgn3430;
        z345_assgn3450 <= z345_assgn345;
        z345_assgn3451 <= z345_assgn3450;
        z80_assgn80 <= z345_assgn3451;
        z349_assgn3490 <= z349_assgn349;
        z82_assgn82 <= z349_assgn3490;
        x3_1_inp_reg <= x3_1_inp;
        r_inp_reg <= r_inp;
        Q1_0_reg <= Q1_0;
        v1_hpc20_reg <= v1_hpc20;
        u0_hpc20_reg <= u0_hpc20;
        p1_hpc20_reg <= p1_hpc20;
        p0_hpc20_reg <= p0_hpc20;
        Q1_1_reg <= Q1_1;
        v0_hpc20_reg <= v0_hpc20;
        u1_hpc20_reg <= u1_hpc20;
        p3_hpc20_reg <= p3_hpc20;
        p2_hpc20_reg <= p2_hpc20;
        L10_0 <= z1_assgn1;
        L10_1 <= z2_assgn2;
        z391_assgn3910 <= z391_assgn391;
        a0_neg_hpc21 <= z391_assgn3910;
        z395_assgn3950 <= z395_assgn395;
        a1_neg_hpc21 <= z395_assgn3950;
        z397_assgn3970 <= z397_assgn397;
        z127_assgn127 <= z397_assgn3970;
        z401_assgn4010 <= z401_assgn401;
        z129_assgn129 <= z401_assgn4010;
        z409_assgn4090 <= z409_assgn409;
        z136_assgn136 <= z409_assgn4090;
        Q4_0_reg <= Q4_0;
        z413_assgn4130 <= z413_assgn413;
        z138_assgn138 <= z413_assgn4130;
        v1_hpc21_reg <= v1_hpc21;
        u0_hpc21_reg <= u0_hpc21;
        p1_hpc21_reg <= p1_hpc21;
        p0_hpc21_reg <= p0_hpc21;
        z421_assgn4210 <= z421_assgn421;
        z144_assgn144 <= z421_assgn4210;
        Q4_1_reg <= Q4_1;
        z425_assgn4250 <= z425_assgn425;
        z146_assgn146 <= z425_assgn4250;
        v0_hpc21_reg <= v0_hpc21;
        u1_hpc21_reg <= u1_hpc21;
        p3_hpc21_reg <= p3_hpc21;
        p2_hpc21_reg <= p2_hpc21;
        T0_0_reg <= T0_0;
        T0_1_reg <= T0_1;
        z453_assgn4530 <= z453_assgn453;
        z453_assgn4531 <= z453_assgn4530;
        z171_assgn171 <= z453_assgn4531;
        z457_assgn4570 <= z457_assgn457;
        z457_assgn4571 <= z457_assgn4570;
        z173_assgn173 <= z457_assgn4571;
        z461_assgn4610 <= z461_assgn461;
        z175_assgn175 <= z461_assgn4610;
        z465_assgn4650 <= z465_assgn465;
        z177_assgn177 <= z465_assgn4650;
        Q3_0_reg <= Q3_0;
        v1_hpc22_reg <= v1_hpc22;
        u0_hpc22_reg <= u0_hpc22;
        p1_hpc22_reg <= p1_hpc22;
        p0_hpc22_reg <= p0_hpc22;
        Q3_1_reg <= Q3_1;
        v0_hpc22_reg <= v0_hpc22;
        u1_hpc22_reg <= u1_hpc22;
        p3_hpc22_reg <= p3_hpc22;
        p2_hpc22_reg <= p2_hpc22;
        z489_assgn4890 <= z489_assgn489;
        z489_assgn4891 <= z489_assgn4890;
        z199_assgn199 <= z489_assgn4891;
        z493_assgn4930 <= z493_assgn493;
        z493_assgn4931 <= z493_assgn4930;
        z201_assgn201 <= z493_assgn4931;
        z497_assgn4970 <= z497_assgn497;
        z203_assgn203 <= z497_assgn4970;
        z501_assgn5010 <= z501_assgn501;
        z205_assgn205 <= z501_assgn5010;
        Q7_0_reg <= Q7_0;
        v1_hpc23_reg <= v1_hpc23;
        u0_hpc23_reg <= u0_hpc23;
        p1_hpc23_reg <= p1_hpc23;
        p0_hpc23_reg <= p0_hpc23;
        Q7_1_reg <= Q7_1;
        v0_hpc23_reg <= v0_hpc23;
        u1_hpc23_reg <= u1_hpc23;
        p3_hpc23_reg <= p3_hpc23;
        p2_hpc23_reg <= p2_hpc23;
        z521_assgn5210 <= z521_assgn521;
        z224_assgn224 <= z521_assgn5210;
        z527_assgn5270 <= z527_assgn527;
        z228_assgn228 <= z527_assgn5270;
        T2_0_reg <= T2_0;
        T2_1_reg <= T2_1;
        z541_assgn5410 <= z541_assgn541;
        z240_assgn240 <= z541_assgn5410;
        Y0_0 <= z9_assgn9;
        Y1_0 <= (L7_0 ^ Y1_01);
        Y2_0 <= z11_assgn11;
        z553_assgn5530 <= z553_assgn553;
        z249_assgn249 <= z553_assgn5530;
        Y3_0 <= z13_assgn13;
        z559_assgn5590 <= z559_assgn559;
        z254_assgn254 <= z559_assgn5590;
        Y0_1 <= z15_assgn15;
        Y1_1 <= (L7_1 ^ Y1_11);
        Y2_1 <= z17_assgn17;
        z571_assgn5710 <= z571_assgn571;
        z263_assgn263 <= z571_assgn5710;
        Y3_1 <= z19_assgn19;
    end

endmodule

