module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r1,
    r2,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r1;
    input  r2;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    reg z3_assgn3;
    wire z243_assgn243;
    reg z243_assgn2430;
    reg x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    reg z5_assgn5;
    wire z253_assgn253;
    reg z253_assgn2530;
    reg x3_1_inp;
    wire r1_inp;
    wire r2_inp;
    reg z7_assgn7;
    reg x1_0_inp_reg;
    wire L0_0;
    wire L1_0;
    wire z265_assgn265;
    reg z265_assgn2650;
    reg z265_assgn2651;
    reg z265_assgn2652;
    reg z51_assgn51;
    wire z267_assgn267;
    reg z267_assgn2670;
    reg z267_assgn2671;
    reg z52_assgn52;
    wire L8_0;
    wire z271_assgn271;
    reg z271_assgn2710;
    reg z54_assgn54;
    wire L5_0;
    reg x1_1_inp_reg;
    wire L0_1;
    wire L1_1;
    wire z279_assgn279;
    reg z279_assgn2790;
    reg z279_assgn2791;
    reg z279_assgn2792;
    reg z59_assgn59;
    wire z281_assgn281;
    reg z281_assgn2810;
    reg z281_assgn2811;
    reg z60_assgn60;
    wire L8_1;
    wire z285_assgn285;
    reg z285_assgn2850;
    reg z62_assgn62;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire z305_assgn305;
    reg z305_assgn3050;
    reg z79_assgn79;
    wire z307_assgn307;
    reg z307_assgn3070;
    reg z307_assgn3071;
    reg z80_assgn80;
    wire L2_0;
    wire z311_assgn311;
    reg z311_assgn3110;
    reg z82_assgn82;
    reg x3_0_inp_reg;
    wire L3_0;
    wire z315_assgn315;
    reg z315_assgn3150;
    reg z83_assgn83;
    wire z317_assgn317;
    reg z317_assgn3170;
    reg z317_assgn3171;
    reg z84_assgn84;
    wire L2_1;
    wire z321_assgn321;
    reg z321_assgn3210;
    reg z86_assgn86;
    reg x3_1_inp_reg;
    wire L3_1;
    wire b0_preshared_hpc10;
    wire b1_preshared_hpc10;
    reg b1_preshared_hpc10_reg;
    wire p2_hpc10;
    wire i1_hpc10;
    reg b0_preshared_hpc10_reg;
    wire p3_hpc10;
    wire i2_hpc10;
    wire z337_assgn337;
    reg z337_assgn3370;
    reg z99_assgn99;
    reg Q0_0_reg;
    wire p1_hpc10;
    wire z341_assgn341;
    reg z341_assgn3410;
    reg z101_assgn101;
    reg Q0_1_reg;
    wire p4_hpc10;
    reg i1_hpc10_reg;
    wire T0_0;
    reg i2_hpc10_reg;
    wire T0_1;
    wire z1_assgn1;
    reg L10_0;
    wire z2_assgn2;
    reg L10_1;
    reg r1_inp_reg;
    wire b0_preshared_hpc11;
    wire b1_preshared_hpc11;
    wire z361_assgn361;
    reg z361_assgn3610;
    reg z120_assgn120;
    reg b1_preshared_hpc11_reg;
    wire p2_hpc11;
    reg z7_assgn7_reg;
    wire i1_hpc11;
    wire z367_assgn367;
    reg z367_assgn3670;
    reg z124_assgn124;
    reg b0_preshared_hpc11_reg;
    wire p3_hpc11;
    wire i2_hpc11;
    wire z373_assgn373;
    reg z373_assgn3730;
    reg z127_assgn127;
    wire z375_assgn375;
    reg z375_assgn3750;
    reg z375_assgn3751;
    reg z128_assgn128;
    wire p1_hpc11;
    wire z379_assgn379;
    reg z379_assgn3790;
    reg z129_assgn129;
    wire z381_assgn381;
    reg z381_assgn3810;
    reg z381_assgn3811;
    reg z130_assgn130;
    wire p4_hpc11;
    reg i1_hpc11_reg;
    wire T2_0;
    reg i2_hpc11_reg;
    wire T2_1;
    reg T0_0_reg;
    wire Q2_0;
    wire L4_0;
    wire Q7_0;
    wire Q6_0;
    reg T0_1_reg;
    wire Q2_1;
    wire L4_1;
    wire Q7_1;
    wire Q6_1;
    wire z405_assgn405;
    reg z405_assgn4050;
    reg z151_assgn151;
    wire b0_preshared_hpc12;
    wire z409_assgn409;
    reg z409_assgn4090;
    reg z153_assgn153;
    wire b1_preshared_hpc12;
    reg b1_preshared_hpc12_reg;
    wire p2_hpc12;
    wire z415_assgn415;
    reg z415_assgn4150;
    reg z157_assgn157;
    wire i1_hpc12;
    reg b0_preshared_hpc12_reg;
    wire p3_hpc12;
    wire z421_assgn421;
    reg z421_assgn4210;
    reg z161_assgn161;
    wire i2_hpc12;
    wire z425_assgn425;
    reg z425_assgn4250;
    reg z163_assgn163;
    reg Q2_0_reg;
    wire p1_hpc12;
    wire z429_assgn429;
    reg z429_assgn4290;
    reg z165_assgn165;
    reg Q2_1_reg;
    wire p4_hpc12;
    reg i1_hpc12_reg;
    wire T1_0;
    reg i2_hpc12_reg;
    wire T1_1;
    wire z437_assgn437;
    reg z437_assgn4370;
    reg z171_assgn171;
    wire b0_preshared_hpc13;
    wire z441_assgn441;
    reg z441_assgn4410;
    reg z173_assgn173;
    wire b1_preshared_hpc13;
    reg b1_preshared_hpc13_reg;
    wire p2_hpc13;
    wire z447_assgn447;
    reg z447_assgn4470;
    reg z177_assgn177;
    wire i1_hpc13;
    reg b0_preshared_hpc13_reg;
    wire p3_hpc13;
    wire z453_assgn453;
    reg z453_assgn4530;
    reg z181_assgn181;
    wire i2_hpc13;
    wire z457_assgn457;
    reg z457_assgn4570;
    reg z183_assgn183;
    reg Q6_0_reg;
    wire p1_hpc13;
    wire z461_assgn461;
    reg z461_assgn4610;
    reg z185_assgn185;
    reg Q6_1_reg;
    wire p4_hpc13;
    reg i1_hpc13_reg;
    wire T3_0;
    reg i2_hpc13_reg;
    wire T3_1;
    wire z469_assgn469;
    reg z469_assgn4690;
    reg z192_assgn192;
    wire L7_0;
    wire L11_0;
    wire z475_assgn475;
    reg z475_assgn4750;
    reg z196_assgn196;
    wire L7_1;
    wire L11_1;
    reg T2_0_reg;
    wire Y0_01;
    wire Y1_01;
    reg T2_1_reg;
    wire Y0_11;
    wire Y1_11;
    wire z489_assgn489;
    reg z489_assgn4890;
    reg z208_assgn208;
    wire z9_assgn9;
    wire z11_assgn11;
    wire z501_assgn501;
    reg z501_assgn5010;
    reg z217_assgn217;
    wire z13_assgn13;
    wire z507_assgn507;
    reg z507_assgn5070;
    reg z222_assgn222;
    wire z15_assgn15;
    wire z17_assgn17;
    wire z519_assgn519;
    reg z519_assgn5190;
    reg z231_assgn231;
    wire z19_assgn19;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign z243_assgn243 = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign z253_assgn253 = x3_1;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign L0_0 = (x1_0_inp_reg ^ z3_assgn3);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign z265_assgn265 = x0_0_inp;
    assign z267_assgn267 = z3_assgn3;
    assign L8_0 = (z52_assgn52 ^ z51_assgn51);
    assign z271_assgn271 = x0_0_inp;
    assign L5_0 = (z54_assgn54 ^ x3_0_inp);
    assign L0_1 = (x1_1_inp_reg ^ z5_assgn5);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign z279_assgn279 = x0_1_inp;
    assign z281_assgn281 = z5_assgn5;
    assign L8_1 = (z60_assgn60 ^ z59_assgn59);
    assign z285_assgn285 = x0_1_inp;
    assign L5_1 = (z62_assgn62 ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !z3_assgn3;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !z5_assgn5;
    assign z305_assgn305 = z3_assgn3;
    assign z307_assgn307 = Q1_0;
    assign L2_0 = (z80_assgn80 ^ z79_assgn79);
    assign z311_assgn311 = Q0_0;
    assign L3_0 = (z82_assgn82 ^ x3_0_inp_reg);
    assign z315_assgn315 = z5_assgn5;
    assign z317_assgn317 = Q1_1;
    assign L2_1 = (z84_assgn84 ^ z83_assgn83);
    assign z321_assgn321 = Q0_1;
    assign L3_1 = (z86_assgn86 ^ x3_1_inp_reg);
    assign b0_preshared_hpc10 = (Q1_0 ^ r1_inp);
    assign b1_preshared_hpc10 = (Q1_1 ^ r1_inp);
    assign p2_hpc10 = (Q0_0 & b1_preshared_hpc10_reg);
    assign i1_hpc10 = (p2_hpc10 ^ z7_assgn7);
    assign p3_hpc10 = (Q0_1 & b0_preshared_hpc10_reg);
    assign i2_hpc10 = (p3_hpc10 ^ z7_assgn7);
    assign z337_assgn337 = b0_preshared_hpc10;
    assign p1_hpc10 = (Q0_0_reg & z99_assgn99);
    assign z341_assgn341 = b1_preshared_hpc10;
    assign p4_hpc10 = (Q0_1_reg & z101_assgn101);
    assign T0_0 = (i1_hpc10_reg ^ p1_hpc10);
    assign T0_1 = (i2_hpc10_reg ^ p4_hpc10);
    assign z1_assgn1 = !L2_0;
    assign z2_assgn2 = !L2_1;
    assign b0_preshared_hpc11 = (Q4_0 ^ r1_inp_reg);
    assign b1_preshared_hpc11 = (Q4_1 ^ r1_inp_reg);
    assign z361_assgn361 = x1_0_inp;
    assign p2_hpc11 = (z120_assgn120 & b1_preshared_hpc11_reg);
    assign i1_hpc11 = (p2_hpc11 ^ z7_assgn7_reg);
    assign z367_assgn367 = x1_1_inp;
    assign p3_hpc11 = (z124_assgn124 & b0_preshared_hpc11_reg);
    assign i2_hpc11 = (p3_hpc11 ^ z7_assgn7_reg);
    assign z373_assgn373 = b0_preshared_hpc11;
    assign z375_assgn375 = x1_0_inp;
    assign p1_hpc11 = (z128_assgn128 & z127_assgn127);
    assign z379_assgn379 = b1_preshared_hpc11;
    assign z381_assgn381 = x1_1_inp;
    assign p4_hpc11 = (z130_assgn130 & z129_assgn129);
    assign T2_0 = (i1_hpc11_reg ^ p1_hpc11);
    assign T2_1 = (i2_hpc11_reg ^ p4_hpc11);
    assign Q2_0 = (T0_0_reg ^ L2_0);
    assign L4_0 = (T0_0_reg ^ T2_0);
    assign Q7_0 = (T0_0 ^ L5_0);
    assign Q6_0 = (L4_0 ^ L3_0);
    assign Q2_1 = (T0_1_reg ^ L2_1);
    assign L4_1 = (T0_1_reg ^ T2_1);
    assign Q7_1 = (T0_1 ^ L5_1);
    assign Q6_1 = (L4_1 ^ L3_1);
    assign z405_assgn405 = r1_inp;
    assign b0_preshared_hpc12 = (Q3_0 ^ z151_assgn151);
    assign z409_assgn409 = r1_inp;
    assign b1_preshared_hpc12 = (Q3_1 ^ z153_assgn153);
    assign p2_hpc12 = (Q2_0 & b1_preshared_hpc12_reg);
    assign z415_assgn415 = z7_assgn7;
    assign i1_hpc12 = (p2_hpc12 ^ z157_assgn157);
    assign p3_hpc12 = (Q2_1 & b0_preshared_hpc12_reg);
    assign z421_assgn421 = z7_assgn7;
    assign i2_hpc12 = (p3_hpc12 ^ z161_assgn161);
    assign z425_assgn425 = b0_preshared_hpc12;
    assign p1_hpc12 = (Q2_0_reg & z163_assgn163);
    assign z429_assgn429 = b1_preshared_hpc12;
    assign p4_hpc12 = (Q2_1_reg & z165_assgn165);
    assign T1_0 = (i1_hpc12_reg ^ p1_hpc12);
    assign T1_1 = (i2_hpc12_reg ^ p4_hpc12);
    assign z437_assgn437 = r1_inp;
    assign b0_preshared_hpc13 = (Q7_0 ^ z171_assgn171);
    assign z441_assgn441 = r1_inp;
    assign b1_preshared_hpc13 = (Q7_1 ^ z173_assgn173);
    assign p2_hpc13 = (Q6_0 & b1_preshared_hpc13_reg);
    assign z447_assgn447 = z7_assgn7;
    assign i1_hpc13 = (p2_hpc13 ^ z177_assgn177);
    assign p3_hpc13 = (Q6_1 & b0_preshared_hpc13_reg);
    assign z453_assgn453 = z7_assgn7;
    assign i2_hpc13 = (p3_hpc13 ^ z181_assgn181);
    assign z457_assgn457 = b0_preshared_hpc13;
    assign p1_hpc13 = (Q6_0_reg & z183_assgn183);
    assign z461_assgn461 = b1_preshared_hpc13;
    assign p4_hpc13 = (Q6_1_reg & z185_assgn185);
    assign T3_0 = (i1_hpc13_reg ^ p1_hpc13);
    assign T3_1 = (i2_hpc13_reg ^ p4_hpc13);
    assign z469_assgn469 = T0_0;
    assign L7_0 = (z192_assgn192 ^ T1_0);
    assign L11_0 = (T1_0 ^ L10_0);
    assign z475_assgn475 = T0_1;
    assign L7_1 = (z196_assgn196 ^ T1_1);
    assign L11_1 = (T1_1 ^ L10_1);
    assign Y0_01 = (L7_0 ^ T2_0_reg);
    assign Y1_01 = (L8_0 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1_reg);
    assign Y1_11 = (L8_1 ^ T3_1);
    assign z489_assgn489 = x3_0_inp;
    assign z9_assgn9 = (z208_assgn208 ^ Y0_01);
    assign z11_assgn11 = (L11_0 ^ T2_0_reg);
    assign z501_assgn501 = L5_0;
    assign z13_assgn13 = (T2_0_reg ^ z217_assgn217);
    assign z507_assgn507 = x3_1_inp;
    assign z15_assgn15 = (z222_assgn222 ^ Y0_11);
    assign z17_assgn17 = (L11_1 ^ T2_1_reg);
    assign z519_assgn519 = L5_1;
    assign z19_assgn19 = (T2_1_reg ^ z231_assgn231);

    always @(posedge clk) begin
        z3_assgn3 <= x2_0_inp;
        z243_assgn2430 <= z243_assgn243;
        x3_0_inp <= z243_assgn2430;
        z5_assgn5 <= x2_1_inp;
        z253_assgn2530 <= z253_assgn253;
        x3_1_inp <= z253_assgn2530;
        z7_assgn7 <= r2_inp;
        x1_0_inp_reg <= x1_0_inp;
        z265_assgn2650 <= z265_assgn265;
        z265_assgn2651 <= z265_assgn2650;
        z265_assgn2652 <= z265_assgn2651;
        z51_assgn51 <= z265_assgn2652;
        z267_assgn2670 <= z267_assgn267;
        z267_assgn2671 <= z267_assgn2670;
        z52_assgn52 <= z267_assgn2671;
        z271_assgn2710 <= z271_assgn271;
        z54_assgn54 <= z271_assgn2710;
        x1_1_inp_reg <= x1_1_inp;
        z279_assgn2790 <= z279_assgn279;
        z279_assgn2791 <= z279_assgn2790;
        z279_assgn2792 <= z279_assgn2791;
        z59_assgn59 <= z279_assgn2792;
        z281_assgn2810 <= z281_assgn281;
        z281_assgn2811 <= z281_assgn2810;
        z60_assgn60 <= z281_assgn2811;
        z285_assgn2850 <= z285_assgn285;
        z62_assgn62 <= z285_assgn2850;
        z305_assgn3050 <= z305_assgn305;
        z79_assgn79 <= z305_assgn3050;
        z307_assgn3070 <= z307_assgn307;
        z307_assgn3071 <= z307_assgn3070;
        z80_assgn80 <= z307_assgn3071;
        z311_assgn3110 <= z311_assgn311;
        z82_assgn82 <= z311_assgn3110;
        x3_0_inp_reg <= x3_0_inp;
        z315_assgn3150 <= z315_assgn315;
        z83_assgn83 <= z315_assgn3150;
        z317_assgn3170 <= z317_assgn317;
        z317_assgn3171 <= z317_assgn3170;
        z84_assgn84 <= z317_assgn3171;
        z321_assgn3210 <= z321_assgn321;
        z86_assgn86 <= z321_assgn3210;
        x3_1_inp_reg <= x3_1_inp;
        b1_preshared_hpc10_reg <= b1_preshared_hpc10;
        b0_preshared_hpc10_reg <= b0_preshared_hpc10;
        z337_assgn3370 <= z337_assgn337;
        z99_assgn99 <= z337_assgn3370;
        Q0_0_reg <= Q0_0;
        z341_assgn3410 <= z341_assgn341;
        z101_assgn101 <= z341_assgn3410;
        Q0_1_reg <= Q0_1;
        i1_hpc10_reg <= i1_hpc10;
        i2_hpc10_reg <= i2_hpc10;
        L10_0 <= z1_assgn1;
        L10_1 <= z2_assgn2;
        r1_inp_reg <= r1_inp;
        z361_assgn3610 <= z361_assgn361;
        z120_assgn120 <= z361_assgn3610;
        b1_preshared_hpc11_reg <= b1_preshared_hpc11;
        z7_assgn7_reg <= z7_assgn7;
        z367_assgn3670 <= z367_assgn367;
        z124_assgn124 <= z367_assgn3670;
        b0_preshared_hpc11_reg <= b0_preshared_hpc11;
        z373_assgn3730 <= z373_assgn373;
        z127_assgn127 <= z373_assgn3730;
        z375_assgn3750 <= z375_assgn375;
        z375_assgn3751 <= z375_assgn3750;
        z128_assgn128 <= z375_assgn3751;
        z379_assgn3790 <= z379_assgn379;
        z129_assgn129 <= z379_assgn3790;
        z381_assgn3810 <= z381_assgn381;
        z381_assgn3811 <= z381_assgn3810;
        z130_assgn130 <= z381_assgn3811;
        i1_hpc11_reg <= i1_hpc11;
        i2_hpc11_reg <= i2_hpc11;
        T0_0_reg <= T0_0;
        T0_1_reg <= T0_1;
        z405_assgn4050 <= z405_assgn405;
        z151_assgn151 <= z405_assgn4050;
        z409_assgn4090 <= z409_assgn409;
        z153_assgn153 <= z409_assgn4090;
        b1_preshared_hpc12_reg <= b1_preshared_hpc12;
        z415_assgn4150 <= z415_assgn415;
        z157_assgn157 <= z415_assgn4150;
        b0_preshared_hpc12_reg <= b0_preshared_hpc12;
        z421_assgn4210 <= z421_assgn421;
        z161_assgn161 <= z421_assgn4210;
        z425_assgn4250 <= z425_assgn425;
        z163_assgn163 <= z425_assgn4250;
        Q2_0_reg <= Q2_0;
        z429_assgn4290 <= z429_assgn429;
        z165_assgn165 <= z429_assgn4290;
        Q2_1_reg <= Q2_1;
        i1_hpc12_reg <= i1_hpc12;
        i2_hpc12_reg <= i2_hpc12;
        z437_assgn4370 <= z437_assgn437;
        z171_assgn171 <= z437_assgn4370;
        z441_assgn4410 <= z441_assgn441;
        z173_assgn173 <= z441_assgn4410;
        b1_preshared_hpc13_reg <= b1_preshared_hpc13;
        z447_assgn4470 <= z447_assgn447;
        z177_assgn177 <= z447_assgn4470;
        b0_preshared_hpc13_reg <= b0_preshared_hpc13;
        z453_assgn4530 <= z453_assgn453;
        z181_assgn181 <= z453_assgn4530;
        z457_assgn4570 <= z457_assgn457;
        z183_assgn183 <= z457_assgn4570;
        Q6_0_reg <= Q6_0;
        z461_assgn4610 <= z461_assgn461;
        z185_assgn185 <= z461_assgn4610;
        Q6_1_reg <= Q6_1;
        i1_hpc13_reg <= i1_hpc13;
        i2_hpc13_reg <= i2_hpc13;
        z469_assgn4690 <= z469_assgn469;
        z192_assgn192 <= z469_assgn4690;
        z475_assgn4750 <= z475_assgn475;
        z196_assgn196 <= z475_assgn4750;
        T2_0_reg <= T2_0;
        T2_1_reg <= T2_1;
        z489_assgn4890 <= z489_assgn489;
        z208_assgn208 <= z489_assgn4890;
        Y0_0 <= z9_assgn9;
        Y1_0 <= (L7_0 ^ Y1_01);
        Y2_0 <= z11_assgn11;
        z501_assgn5010 <= z501_assgn501;
        z217_assgn217 <= z501_assgn5010;
        Y3_0 <= z13_assgn13;
        z507_assgn5070 <= z507_assgn507;
        z222_assgn222 <= z507_assgn5070;
        Y0_1 <= z15_assgn15;
        Y1_1 <= (L7_1 ^ Y1_11);
        Y2_1 <= z17_assgn17;
        z519_assgn5190 <= z519_assgn519;
        z231_assgn231 <= z519_assgn5190;
        Y3_1 <= z19_assgn19;
    end

endmodule

