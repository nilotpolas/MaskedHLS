module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r0,
    r1,
    r0_1,
    r1_1,
    r2_1,
    r3_1,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r0;
    input  r1;
    input  r0_1;
    input  r1_1;
    input  r2_1;
    input  r3_1;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    wire x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    wire x3_1_inp;
    wire r0_inp;
    wire r1_inp;
    wire r0_1_inp;
    wire r1_1_inp;
    wire r2_1_inp;
    wire r3_1_inp;
    wire L0_0;
    wire L1_0;
    wire L8_0;
    wire L5_0;
    wire L0_1;
    wire L1_1;
    wire L8_1;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire L2_0;
    wire L3_0;
    wire L2_1;
    wire L3_1;
    wire m0_comar0;
    wire m1_comar0;
    wire m2_comar0;
    wire m3_comar0;
    reg m0_comar0_reg;
    reg m1_comar0_reg;
    wire p2_comar0;
    reg m3_comar0_reg;
    reg m2_comar0_reg;
    wire p3_comar0;
    wire p1_comar0;
    wire p4_comar0;
    reg r0_1_inp_reg;
    wire i0_comar0;
    reg r1_1_inp_reg;
    wire i1_comar0;
    reg r2_1_inp_reg;
    wire i2_comar0;
    reg r3_1_inp_reg;
    wire i3_comar0;
    reg i1_comar0_reg;
    reg i2_comar0_reg;
    wire i1xori2_comar0;
    reg i0_comar0_reg;
    reg i3_comar0_reg;
    wire i0xori3_comar0;
    reg T0_0;
    wire y1_1_comar0;
    wire y1_2_comar0;
    wire y1_3_comar0;
    wire y1_4_comar0;
    wire T0_1;
    wire L10_0;
    wire L10_1;
    wire m0_comar1;
    wire m1_comar1;
    wire m2_comar1;
    wire m3_comar1;
    reg m0_comar1_reg;
    reg m1_comar1_reg;
    wire p2_comar1;
    reg m3_comar1_reg;
    reg m2_comar1_reg;
    wire p3_comar1;
    wire p1_comar1;
    wire p4_comar1;
    wire i0_comar1;
    wire i1_comar1;
    wire i2_comar1;
    wire i3_comar1;
    reg i1_comar1_reg;
    reg i2_comar1_reg;
    wire i1xori2_comar1;
    reg i0_comar1_reg;
    reg i3_comar1_reg;
    wire i0xori3_comar1;
    reg T2_0;
    wire y1_1_comar1;
    wire y1_2_comar1;
    wire y1_3_comar1;
    wire y1_4_comar1;
    wire T2_1;
    wire z445_assgn445;
    reg z445_assgn4450;
    reg z445_assgn4451;
    reg z159_assgn159;
    wire Q2_0;
    wire L4_0;
    wire z451_assgn451;
    reg z451_assgn4510;
    reg z451_assgn4511;
    reg z163_assgn163;
    wire Q7_0;
    wire z455_assgn455;
    reg z455_assgn4550;
    reg z455_assgn4551;
    reg z165_assgn165;
    wire Q6_0;
    wire Q2_1;
    wire L4_1;
    wire Q7_1;
    wire Q6_1;
    wire z467_assgn467;
    reg z467_assgn4670;
    reg z467_assgn4671;
    reg z175_assgn175;
    wire m0_comar2;
    wire m1_comar2;
    wire m2_comar2;
    wire m3_comar2;
    wire z477_assgn477;
    reg z477_assgn4770;
    reg z477_assgn4771;
    reg z477_assgn4772;
    reg z183_assgn183;
    reg m0_comar2_reg;
    wire p2_comar2;
    reg m3_comar2_reg;
    reg m2_comar2_reg;
    wire p3_comar2;
    wire z483_assgn483;
    reg z483_assgn4830;
    reg z483_assgn4831;
    reg z483_assgn4832;
    reg z187_assgn187;
    wire p1_comar2;
    reg m1_comar2_reg;
    wire p4_comar2;
    wire z489_assgn489;
    reg z489_assgn4890;
    reg z489_assgn4891;
    reg z489_assgn4892;
    reg z191_assgn191;
    wire i0_comar2;
    wire z493_assgn493;
    reg z493_assgn4930;
    reg z493_assgn4931;
    reg z493_assgn4932;
    reg z193_assgn193;
    wire i1_comar2;
    wire i2_comar2;
    wire i3_comar2;
    wire z501_assgn501;
    reg z501_assgn5010;
    reg z501_assgn5011;
    reg z501_assgn5012;
    reg z199_assgn199;
    reg i1_comar2_reg;
    wire i1xori2_comar2;
    wire z505_assgn505;
    reg z505_assgn5050;
    reg z505_assgn5051;
    reg z505_assgn5052;
    reg z201_assgn201;
    reg i0_comar2_reg;
    wire i0xori3_comar2;
    reg T1_0;
    wire y1_1_comar2;
    wire y1_2_comar2;
    wire y1_3_comar2;
    wire y1_4_comar2;
    wire T1_1;
    wire z521_assgn521;
    reg z521_assgn5210;
    reg z521_assgn5211;
    reg z215_assgn215;
    wire m0_comar3;
    wire m1_comar3;
    wire z527_assgn527;
    reg z527_assgn5270;
    reg z527_assgn5271;
    reg z219_assgn219;
    wire m2_comar3;
    wire m3_comar3;
    wire z533_assgn533;
    reg z533_assgn5330;
    reg z533_assgn5331;
    reg z533_assgn5332;
    reg z223_assgn223;
    reg m0_comar3_reg;
    wire p2_comar3;
    wire z537_assgn537;
    reg z537_assgn5370;
    reg z537_assgn5371;
    reg z537_assgn5372;
    reg z226_assgn226;
    reg m2_comar3_reg;
    wire p3_comar3;
    wire p1_comar3;
    reg m3_comar3_reg;
    reg m1_comar3_reg;
    wire p4_comar3;
    wire z545_assgn545;
    reg z545_assgn5450;
    reg z545_assgn5451;
    reg z545_assgn5452;
    reg z231_assgn231;
    wire i0_comar3;
    wire z549_assgn549;
    reg z549_assgn5490;
    reg z549_assgn5491;
    reg z549_assgn5492;
    reg z233_assgn233;
    wire i1_comar3;
    wire z553_assgn553;
    reg z553_assgn5530;
    reg z553_assgn5531;
    reg z553_assgn5532;
    reg z235_assgn235;
    wire i2_comar3;
    wire i3_comar3;
    reg i1_comar3_reg;
    reg i2_comar3_reg;
    wire i1xori2_comar3;
    wire z561_assgn561;
    reg z561_assgn5610;
    reg z561_assgn5611;
    reg z561_assgn5612;
    reg z241_assgn241;
    reg i0_comar3_reg;
    wire i0xori3_comar3;
    reg T3_0;
    wire y1_1_comar3;
    wire y1_2_comar3;
    wire y1_3_comar3;
    wire y1_4_comar3;
    wire T3_1;
    wire z577_assgn577;
    reg z577_assgn5770;
    reg z577_assgn5771;
    reg z256_assgn256;
    wire L7_0;
    wire z581_assgn581;
    reg z581_assgn5810;
    reg z581_assgn5811;
    reg z581_assgn5812;
    reg z581_assgn5813;
    reg z581_assgn5814;
    reg z257_assgn257;
    wire L11_0;
    wire L7_1;
    wire L11_1;
    wire z589_assgn589;
    reg z589_assgn5890;
    reg z589_assgn5891;
    reg z263_assgn263;
    wire Y0_01;
    wire z593_assgn593;
    reg z593_assgn5930;
    reg z593_assgn5931;
    reg z593_assgn5932;
    reg z593_assgn5933;
    reg z593_assgn5934;
    reg z266_assgn266;
    wire Y1_01;
    wire Y0_11;
    wire Y1_11;
    wire z601_assgn601;
    reg z601_assgn6010;
    reg z601_assgn6011;
    reg z601_assgn6012;
    reg z601_assgn6013;
    reg z601_assgn6014;
    reg z272_assgn272;
    wire z1_assgn1;
    wire z609_assgn609;
    reg z609_assgn6090;
    reg z609_assgn6091;
    reg z277_assgn277;
    wire z3_assgn3;
    wire z615_assgn615;
    reg z615_assgn6150;
    reg z615_assgn6151;
    reg z281_assgn281;
    wire z5_assgn5;
    wire z619_assgn619;
    reg z619_assgn6190;
    reg z619_assgn6191;
    reg z619_assgn6192;
    wire z621_assgn621;
    reg z621_assgn6210;
    reg z621_assgn6211;
    reg z621_assgn6212;
    reg z621_assgn6213;
    reg z621_assgn6214;
    reg z621_assgn6215;
    wire z623_assgn623;
    reg z623_assgn6230;
    reg z623_assgn6231;
    reg z623_assgn6232;
    reg z623_assgn6233;
    reg z623_assgn6234;
    reg z623_assgn6235;
    wire z625_assgn625;
    reg z625_assgn6250;
    reg z625_assgn6251;
    reg z625_assgn6252;
    reg z625_assgn6253;
    reg z625_assgn6254;
    reg z625_assgn6255;
    wire z627_assgn627;
    reg z627_assgn6270;
    reg z627_assgn6271;
    reg z627_assgn6272;
    reg z627_assgn6273;
    reg z627_assgn6274;
    reg z627_assgn6275;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign x3_0_inp = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign x3_1_inp = x3_1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r0_1_inp = r0_1;
    assign r1_1_inp = r1_1;
    assign r2_1_inp = r2_1;
    assign r3_1_inp = r3_1;
    assign L0_0 = (x1_0_inp ^ x2_0_inp);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign L8_0 = (x2_0_inp ^ x0_0_inp);
    assign L5_0 = (x0_0_inp ^ x3_0_inp);
    assign L0_1 = (x1_1_inp ^ x2_1_inp);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign L8_1 = (x2_1_inp ^ x0_1_inp);
    assign L5_1 = (x0_1_inp ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !x2_0_inp;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !x2_1_inp;
    assign L2_0 = (Q1_0 ^ x2_0_inp);
    assign L3_0 = (Q0_0 ^ x3_0_inp);
    assign L2_1 = (Q1_1 ^ x2_1_inp);
    assign L3_1 = (Q0_1 ^ x3_1_inp);
    assign m0_comar0 = (Q0_0 ^ r0_inp);
    assign m1_comar0 = (Q1_1 ^ r1_inp);
    assign m2_comar0 = (Q1_0 ^ r1_inp);
    assign m3_comar0 = (Q0_1 ^ r0_inp);
    assign p2_comar0 = (m0_comar0_reg & m1_comar0_reg);
    assign p3_comar0 = (m3_comar0_reg & m2_comar0_reg);
    assign p1_comar0 = (m0_comar0_reg & m2_comar0_reg);
    assign p4_comar0 = (m3_comar0_reg & m1_comar0_reg);
    assign i0_comar0 = (p1_comar0 ^ r0_1_inp_reg);
    assign i1_comar0 = (p2_comar0 ^ r1_1_inp_reg);
    assign i2_comar0 = (p3_comar0 ^ r2_1_inp_reg);
    assign i3_comar0 = (p4_comar0 ^ r3_1_inp_reg);
    assign i1xori2_comar0 = (i1_comar0_reg ^ i2_comar0_reg);
    assign i0xori3_comar0 = (i0_comar0_reg ^ i3_comar0_reg);
    assign y1_1_comar0 = (r0_inp ^ r0_inp);
    assign y1_2_comar0 = (y1_1_comar0 ^ r0_1_inp);
    assign y1_3_comar0 = (y1_2_comar0 ^ r1_1_inp);
    assign y1_4_comar0 = (y1_3_comar0 ^ r2_1_inp);
    assign T0_1 = (y1_4_comar0 ^ r3_1_inp);
    assign L10_0 = !L2_0;
    assign L10_1 = !L2_1;
    assign m0_comar1 = (x1_0_inp ^ r0_inp);
    assign m1_comar1 = (Q4_1 ^ r1_inp);
    assign m2_comar1 = (Q4_0 ^ r1_inp);
    assign m3_comar1 = (x1_1_inp ^ r0_inp);
    assign p2_comar1 = (m0_comar1_reg & m1_comar1_reg);
    assign p3_comar1 = (m3_comar1_reg & m2_comar1_reg);
    assign p1_comar1 = (m0_comar1_reg & m2_comar1_reg);
    assign p4_comar1 = (m3_comar1_reg & m1_comar1_reg);
    assign i0_comar1 = (p1_comar1 ^ r0_1_inp_reg);
    assign i1_comar1 = (p2_comar1 ^ r1_1_inp_reg);
    assign i2_comar1 = (p3_comar1 ^ r2_1_inp_reg);
    assign i3_comar1 = (p4_comar1 ^ r3_1_inp_reg);
    assign i1xori2_comar1 = (i1_comar1_reg ^ i2_comar1_reg);
    assign i0xori3_comar1 = (i0_comar1_reg ^ i3_comar1_reg);
    assign y1_1_comar1 = (r0_inp ^ r0_inp);
    assign y1_2_comar1 = (y1_1_comar1 ^ r0_1_inp);
    assign y1_3_comar1 = (y1_2_comar1 ^ r1_1_inp);
    assign y1_4_comar1 = (y1_3_comar1 ^ r2_1_inp);
    assign T2_1 = (y1_4_comar1 ^ r3_1_inp);
    assign z445_assgn445 = L2_0;
    assign Q2_0 = (T0_0 ^ z159_assgn159);
    assign L4_0 = (T0_0 ^ T2_0);
    assign z451_assgn451 = L5_0;
    assign Q7_0 = (T0_0 ^ z163_assgn163);
    assign z455_assgn455 = L3_0;
    assign Q6_0 = (L4_0 ^ z165_assgn165);
    assign Q2_1 = (T0_1 ^ L2_1);
    assign L4_1 = (T0_1 ^ T2_1);
    assign Q7_1 = (T0_1 ^ L5_1);
    assign Q6_1 = (L4_1 ^ L3_1);
    assign z467_assgn467 = r0_inp;
    assign m0_comar2 = (Q2_0 ^ z175_assgn175);
    assign m1_comar2 = (Q3_1 ^ r1_inp);
    assign m2_comar2 = (Q3_0 ^ r1_inp);
    assign m3_comar2 = (Q2_1 ^ r0_inp);
    assign z477_assgn477 = m1_comar2;
    assign p2_comar2 = (m0_comar2_reg & z183_assgn183);
    assign p3_comar2 = (m3_comar2_reg & m2_comar2_reg);
    assign z483_assgn483 = m2_comar2;
    assign p1_comar2 = (m0_comar2_reg & z187_assgn187);
    assign p4_comar2 = (m3_comar2_reg & m1_comar2_reg);
    assign z489_assgn489 = r0_1_inp;
    assign i0_comar2 = (p1_comar2 ^ z191_assgn191);
    assign z493_assgn493 = r1_1_inp;
    assign i1_comar2 = (p2_comar2 ^ z193_assgn193);
    assign i2_comar2 = (p3_comar2 ^ r2_1_inp_reg);
    assign i3_comar2 = (p4_comar2 ^ r3_1_inp_reg);
    assign z501_assgn501 = i2_comar2;
    assign i1xori2_comar2 = (i1_comar2_reg ^ z199_assgn199);
    assign z505_assgn505 = i3_comar2;
    assign i0xori3_comar2 = (i0_comar2_reg ^ z201_assgn201);
    assign y1_1_comar2 = (r0_inp ^ r0_inp);
    assign y1_2_comar2 = (y1_1_comar2 ^ r0_1_inp);
    assign y1_3_comar2 = (y1_2_comar2 ^ r1_1_inp);
    assign y1_4_comar2 = (y1_3_comar2 ^ r2_1_inp);
    assign T1_1 = (y1_4_comar2 ^ r3_1_inp);
    assign z521_assgn521 = r0_inp;
    assign m0_comar3 = (Q6_0 ^ z215_assgn215);
    assign m1_comar3 = (Q7_1 ^ r1_inp);
    assign z527_assgn527 = r1_inp;
    assign m2_comar3 = (Q7_0 ^ z219_assgn219);
    assign m3_comar3 = (Q6_1 ^ r0_inp);
    assign z533_assgn533 = m1_comar3;
    assign p2_comar3 = (m0_comar3_reg & z223_assgn223);
    assign z537_assgn537 = m3_comar3;
    assign p3_comar3 = (z226_assgn226 & m2_comar3_reg);
    assign p1_comar3 = (m0_comar3_reg & m2_comar3_reg);
    assign p4_comar3 = (m3_comar3_reg & m1_comar3_reg);
    assign z545_assgn545 = r0_1_inp;
    assign i0_comar3 = (p1_comar3 ^ z231_assgn231);
    assign z549_assgn549 = r1_1_inp;
    assign i1_comar3 = (p2_comar3 ^ z233_assgn233);
    assign z553_assgn553 = r2_1_inp;
    assign i2_comar3 = (p3_comar3 ^ z235_assgn235);
    assign i3_comar3 = (p4_comar3 ^ r3_1_inp_reg);
    assign i1xori2_comar3 = (i1_comar3_reg ^ i2_comar3_reg);
    assign z561_assgn561 = i3_comar3;
    assign i0xori3_comar3 = (i0_comar3_reg ^ z241_assgn241);
    assign y1_1_comar3 = (r0_inp ^ r0_inp);
    assign y1_2_comar3 = (y1_1_comar3 ^ r0_1_inp);
    assign y1_3_comar3 = (y1_2_comar3 ^ r1_1_inp);
    assign y1_4_comar3 = (y1_3_comar3 ^ r2_1_inp);
    assign T3_1 = (y1_4_comar3 ^ r3_1_inp);
    assign z577_assgn577 = T0_0;
    assign L7_0 = (z256_assgn256 ^ T1_0);
    assign z581_assgn581 = L10_0;
    assign L11_0 = (T1_0 ^ z257_assgn257);
    assign L7_1 = (T0_1 ^ T1_1);
    assign L11_1 = (T1_1 ^ L10_1);
    assign z589_assgn589 = T2_0;
    assign Y0_01 = (L7_0 ^ z263_assgn263);
    assign z593_assgn593 = L8_0;
    assign Y1_01 = (z266_assgn266 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1);
    assign Y1_11 = (L8_1 ^ T3_1);
    assign z601_assgn601 = x3_0_inp;
    assign z1_assgn1 = (z272_assgn272 ^ Y0_01);
    assign z609_assgn609 = T2_0;
    assign z3_assgn3 = (L11_0 ^ z277_assgn277);
    assign z615_assgn615 = L5_0;
    assign z5_assgn5 = (T2_0 ^ z281_assgn281);
    assign z619_assgn619 = z5_assgn5;
    assign z621_assgn621 = (x3_1_inp ^ Y0_11);
    assign z623_assgn623 = (L7_1 ^ Y1_11);
    assign z625_assgn625 = (L11_1 ^ T2_1);
    assign z627_assgn627 = (T2_1 ^ L5_1);

    always @(posedge clk) begin
        m0_comar0_reg <= m0_comar0;
        m1_comar0_reg <= m1_comar0;
        m3_comar0_reg <= m3_comar0;
        m2_comar0_reg <= m2_comar0;
        r0_1_inp_reg <= r0_1_inp;
        r1_1_inp_reg <= r1_1_inp;
        r2_1_inp_reg <= r2_1_inp;
        r3_1_inp_reg <= r3_1_inp;
        i1_comar0_reg <= i1_comar0;
        i2_comar0_reg <= i2_comar0;
        i0_comar0_reg <= i0_comar0;
        i3_comar0_reg <= i3_comar0;
        T0_0 <= (i1xori2_comar0 ^ i0xori3_comar0);
        m0_comar1_reg <= m0_comar1;
        m1_comar1_reg <= m1_comar1;
        m3_comar1_reg <= m3_comar1;
        m2_comar1_reg <= m2_comar1;
        i1_comar1_reg <= i1_comar1;
        i2_comar1_reg <= i2_comar1;
        i0_comar1_reg <= i0_comar1;
        i3_comar1_reg <= i3_comar1;
        T2_0 <= (i1xori2_comar1 ^ i0xori3_comar1);
        z445_assgn4450 <= z445_assgn445;
        z445_assgn4451 <= z445_assgn4450;
        z159_assgn159 <= z445_assgn4451;
        z451_assgn4510 <= z451_assgn451;
        z451_assgn4511 <= z451_assgn4510;
        z163_assgn163 <= z451_assgn4511;
        z455_assgn4550 <= z455_assgn455;
        z455_assgn4551 <= z455_assgn4550;
        z165_assgn165 <= z455_assgn4551;
        z467_assgn4670 <= z467_assgn467;
        z467_assgn4671 <= z467_assgn4670;
        z175_assgn175 <= z467_assgn4671;
        z477_assgn4770 <= z477_assgn477;
        z477_assgn4771 <= z477_assgn4770;
        z477_assgn4772 <= z477_assgn4771;
        z183_assgn183 <= z477_assgn4772;
        m0_comar2_reg <= m0_comar2;
        m3_comar2_reg <= m3_comar2;
        m2_comar2_reg <= m2_comar2;
        z483_assgn4830 <= z483_assgn483;
        z483_assgn4831 <= z483_assgn4830;
        z483_assgn4832 <= z483_assgn4831;
        z187_assgn187 <= z483_assgn4832;
        m1_comar2_reg <= m1_comar2;
        z489_assgn4890 <= z489_assgn489;
        z489_assgn4891 <= z489_assgn4890;
        z489_assgn4892 <= z489_assgn4891;
        z191_assgn191 <= z489_assgn4892;
        z493_assgn4930 <= z493_assgn493;
        z493_assgn4931 <= z493_assgn4930;
        z493_assgn4932 <= z493_assgn4931;
        z193_assgn193 <= z493_assgn4932;
        z501_assgn5010 <= z501_assgn501;
        z501_assgn5011 <= z501_assgn5010;
        z501_assgn5012 <= z501_assgn5011;
        z199_assgn199 <= z501_assgn5012;
        i1_comar2_reg <= i1_comar2;
        z505_assgn5050 <= z505_assgn505;
        z505_assgn5051 <= z505_assgn5050;
        z505_assgn5052 <= z505_assgn5051;
        z201_assgn201 <= z505_assgn5052;
        i0_comar2_reg <= i0_comar2;
        T1_0 <= (i1xori2_comar2 ^ i0xori3_comar2);
        z521_assgn5210 <= z521_assgn521;
        z521_assgn5211 <= z521_assgn5210;
        z215_assgn215 <= z521_assgn5211;
        z527_assgn5270 <= z527_assgn527;
        z527_assgn5271 <= z527_assgn5270;
        z219_assgn219 <= z527_assgn5271;
        z533_assgn5330 <= z533_assgn533;
        z533_assgn5331 <= z533_assgn5330;
        z533_assgn5332 <= z533_assgn5331;
        z223_assgn223 <= z533_assgn5332;
        m0_comar3_reg <= m0_comar3;
        z537_assgn5370 <= z537_assgn537;
        z537_assgn5371 <= z537_assgn5370;
        z537_assgn5372 <= z537_assgn5371;
        z226_assgn226 <= z537_assgn5372;
        m2_comar3_reg <= m2_comar3;
        m3_comar3_reg <= m3_comar3;
        m1_comar3_reg <= m1_comar3;
        z545_assgn5450 <= z545_assgn545;
        z545_assgn5451 <= z545_assgn5450;
        z545_assgn5452 <= z545_assgn5451;
        z231_assgn231 <= z545_assgn5452;
        z549_assgn5490 <= z549_assgn549;
        z549_assgn5491 <= z549_assgn5490;
        z549_assgn5492 <= z549_assgn5491;
        z233_assgn233 <= z549_assgn5492;
        z553_assgn5530 <= z553_assgn553;
        z553_assgn5531 <= z553_assgn5530;
        z553_assgn5532 <= z553_assgn5531;
        z235_assgn235 <= z553_assgn5532;
        i1_comar3_reg <= i1_comar3;
        i2_comar3_reg <= i2_comar3;
        z561_assgn5610 <= z561_assgn561;
        z561_assgn5611 <= z561_assgn5610;
        z561_assgn5612 <= z561_assgn5611;
        z241_assgn241 <= z561_assgn5612;
        i0_comar3_reg <= i0_comar3;
        T3_0 <= (i1xori2_comar3 ^ i0xori3_comar3);
        z577_assgn5770 <= z577_assgn577;
        z577_assgn5771 <= z577_assgn5770;
        z256_assgn256 <= z577_assgn5771;
        z581_assgn5810 <= z581_assgn581;
        z581_assgn5811 <= z581_assgn5810;
        z581_assgn5812 <= z581_assgn5811;
        z581_assgn5813 <= z581_assgn5812;
        z581_assgn5814 <= z581_assgn5813;
        z257_assgn257 <= z581_assgn5814;
        z589_assgn5890 <= z589_assgn589;
        z589_assgn5891 <= z589_assgn5890;
        z263_assgn263 <= z589_assgn5891;
        z593_assgn5930 <= z593_assgn593;
        z593_assgn5931 <= z593_assgn5930;
        z593_assgn5932 <= z593_assgn5931;
        z593_assgn5933 <= z593_assgn5932;
        z593_assgn5934 <= z593_assgn5933;
        z266_assgn266 <= z593_assgn5934;
        z601_assgn6010 <= z601_assgn601;
        z601_assgn6011 <= z601_assgn6010;
        z601_assgn6012 <= z601_assgn6011;
        z601_assgn6013 <= z601_assgn6012;
        z601_assgn6014 <= z601_assgn6013;
        z272_assgn272 <= z601_assgn6014;
        Y0_0 <= z1_assgn1;
        Y1_0 <= (L7_0 ^ Y1_01);
        z609_assgn6090 <= z609_assgn609;
        z609_assgn6091 <= z609_assgn6090;
        z277_assgn277 <= z609_assgn6091;
        Y2_0 <= z3_assgn3;
        z615_assgn6150 <= z615_assgn615;
        z615_assgn6151 <= z615_assgn6150;
        z281_assgn281 <= z615_assgn6151;
        z619_assgn6190 <= z619_assgn619;
        z619_assgn6191 <= z619_assgn6190;
        z619_assgn6192 <= z619_assgn6191;
        Y3_0 <= z619_assgn6192;
        z621_assgn6210 <= z621_assgn621;
        z621_assgn6211 <= z621_assgn6210;
        z621_assgn6212 <= z621_assgn6211;
        z621_assgn6213 <= z621_assgn6212;
        z621_assgn6214 <= z621_assgn6213;
        z621_assgn6215 <= z621_assgn6214;
        Y0_1 <= z621_assgn6215;
        z623_assgn6230 <= z623_assgn623;
        z623_assgn6231 <= z623_assgn6230;
        z623_assgn6232 <= z623_assgn6231;
        z623_assgn6233 <= z623_assgn6232;
        z623_assgn6234 <= z623_assgn6233;
        z623_assgn6235 <= z623_assgn6234;
        Y1_1 <= z623_assgn6235;
        z625_assgn6250 <= z625_assgn625;
        z625_assgn6251 <= z625_assgn6250;
        z625_assgn6252 <= z625_assgn6251;
        z625_assgn6253 <= z625_assgn6252;
        z625_assgn6254 <= z625_assgn6253;
        z625_assgn6255 <= z625_assgn6254;
        Y2_1 <= z625_assgn6255;
        z627_assgn6270 <= z627_assgn627;
        z627_assgn6271 <= z627_assgn6270;
        z627_assgn6272 <= z627_assgn6271;
        z627_assgn6273 <= z627_assgn6272;
        z627_assgn6274 <= z627_assgn6273;
        z627_assgn6275 <= z627_assgn6274;
        Y3_1 <= z627_assgn6275;
    end

endmodule

