module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r1,
    r2,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r1;
    input  r2;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    wire x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    wire x3_1_inp;
    wire r1_inp;
    wire r2_inp;
    wire L0_0;
    wire L1_0;
    wire L8_0;
    wire L5_0;
    wire L0_1;
    wire L1_1;
    wire L8_1;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire L2_0;
    wire L3_0;
    wire L2_1;
    wire L3_1;
    wire b0_preshared_hpc10;
    wire b1_preshared_hpc10;
    reg Q0_0_reg;
    reg b1_preshared_hpc10_reg;
    wire p2_hpc10;
    reg r2_inp_reg;
    wire i1_hpc10;
    reg Q0_1_reg;
    reg b0_preshared_hpc10_reg;
    wire p3_hpc10;
    wire i2_hpc10;
    wire p1_hpc10;
    wire p4_hpc10;
    reg i1_hpc10_reg;
    reg p1_hpc10_reg;
    wire T0_0;
    reg i2_hpc10_reg;
    reg p4_hpc10_reg;
    wire T0_1;
    wire L10_0;
    wire L10_1;
    wire b0_preshared_hpc11;
    wire b1_preshared_hpc11;
    reg x1_0_inp_reg;
    reg b1_preshared_hpc11_reg;
    wire p2_hpc11;
    wire i1_hpc11;
    reg x1_1_inp_reg;
    reg b0_preshared_hpc11_reg;
    wire p3_hpc11;
    wire i2_hpc11;
    wire p1_hpc11;
    wire p4_hpc11;
    reg i1_hpc11_reg;
    reg p1_hpc11_reg;
    wire T2_0;
    reg i2_hpc11_reg;
    reg p4_hpc11_reg;
    wire T2_1;
    wire z329_assgn329;
    reg z329_assgn3290;
    reg z121_assgn121;
    wire Q2_0;
    wire L4_0;
    wire z335_assgn335;
    reg z335_assgn3350;
    reg z125_assgn125;
    wire Q7_0;
    wire z339_assgn339;
    reg z339_assgn3390;
    reg z127_assgn127;
    wire Q6_0;
    wire z343_assgn343;
    reg z343_assgn3430;
    reg z129_assgn129;
    wire Q2_1;
    wire L4_1;
    wire z349_assgn349;
    reg z349_assgn3490;
    reg z133_assgn133;
    wire Q7_1;
    wire z353_assgn353;
    reg z353_assgn3530;
    reg z135_assgn135;
    wire Q6_1;
    wire b0_preshared_hpc12;
    wire b1_preshared_hpc12;
    wire z361_assgn361;
    reg z361_assgn3610;
    reg z141_assgn141;
    wire p2_hpc12;
    wire z365_assgn365;
    reg z365_assgn3650;
    reg z143_assgn143;
    wire i1_hpc12;
    wire z369_assgn369;
    reg z369_assgn3690;
    reg z145_assgn145;
    wire p3_hpc12;
    wire z373_assgn373;
    reg z373_assgn3730;
    reg z147_assgn147;
    wire i2_hpc12;
    wire z377_assgn377;
    reg z377_assgn3770;
    reg z149_assgn149;
    wire p1_hpc12;
    wire z381_assgn381;
    reg z381_assgn3810;
    reg z151_assgn151;
    wire p4_hpc12;
    reg i1_hpc12_reg;
    reg p1_hpc12_reg;
    wire T1_0;
    reg i2_hpc12_reg;
    reg p4_hpc12_reg;
    wire T1_1;
    wire z389_assgn389;
    reg z389_assgn3890;
    reg z157_assgn157;
    wire b0_preshared_hpc13;
    wire z393_assgn393;
    reg z393_assgn3930;
    reg z159_assgn159;
    wire b1_preshared_hpc13;
    reg Q6_0_reg;
    reg b1_preshared_hpc13_reg;
    wire p2_hpc13;
    wire z399_assgn399;
    reg z399_assgn3990;
    reg z399_assgn3991;
    reg z163_assgn163;
    wire i1_hpc13;
    reg Q6_1_reg;
    reg b0_preshared_hpc13_reg;
    wire p3_hpc13;
    wire z405_assgn405;
    reg z405_assgn4050;
    reg z405_assgn4051;
    reg z167_assgn167;
    wire i2_hpc13;
    wire p1_hpc13;
    wire p4_hpc13;
    reg i1_hpc13_reg;
    reg p1_hpc13_reg;
    wire T3_0;
    reg i2_hpc13_reg;
    reg p4_hpc13_reg;
    wire T3_1;
    reg T0_0_reg;
    wire L7_0;
    wire z419_assgn419;
    reg z419_assgn4190;
    reg z419_assgn4191;
    reg z179_assgn179;
    wire L11_0;
    reg T0_1_reg;
    wire L7_1;
    wire z425_assgn425;
    reg z425_assgn4250;
    reg z425_assgn4251;
    reg z183_assgn183;
    wire L11_1;
    reg T2_0_reg;
    wire Y0_01;
    wire z431_assgn431;
    reg z431_assgn4310;
    reg z431_assgn4311;
    reg z431_assgn4312;
    reg z188_assgn188;
    wire Y1_01;
    reg T2_1_reg;
    wire Y0_11;
    wire z437_assgn437;
    reg z437_assgn4370;
    reg z437_assgn4371;
    reg z437_assgn4372;
    reg z192_assgn192;
    wire Y1_11;
    wire z441_assgn441;
    reg z441_assgn4410;
    reg z441_assgn4411;
    reg z194_assgn194;
    wire z1_assgn1;
    wire z445_assgn445;
    reg z445_assgn4450;
    reg L7_0_reg;
    wire z3_assgn3;
    wire z5_assgn5;
    wire z453_assgn453;
    reg z453_assgn4530;
    wire z455_assgn455;
    reg z455_assgn4550;
    reg z205_assgn205;
    wire z7_assgn7;
    wire z459_assgn459;
    reg z459_assgn4590;
    reg z459_assgn4591;
    wire z461_assgn461;
    reg z461_assgn4610;
    reg z461_assgn4611;
    reg z210_assgn210;
    wire z9_assgn9;
    wire z465_assgn465;
    reg z465_assgn4650;
    reg L7_1_reg;
    wire z11_assgn11;
    wire z13_assgn13;
    wire z473_assgn473;
    reg z473_assgn4730;
    wire z475_assgn475;
    reg z475_assgn4750;
    reg z221_assgn221;
    wire z15_assgn15;
    wire z479_assgn479;
    reg z479_assgn4790;
    reg z479_assgn4791;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign x3_0_inp = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign x3_1_inp = x3_1;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign L0_0 = (x1_0_inp ^ x2_0_inp);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign L8_0 = (x2_0_inp ^ x0_0_inp);
    assign L5_0 = (x0_0_inp ^ x3_0_inp);
    assign L0_1 = (x1_1_inp ^ x2_1_inp);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign L8_1 = (x2_1_inp ^ x0_1_inp);
    assign L5_1 = (x0_1_inp ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !x2_0_inp;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !x2_1_inp;
    assign L2_0 = (Q1_0 ^ x2_0_inp);
    assign L3_0 = (Q0_0 ^ x3_0_inp);
    assign L2_1 = (Q1_1 ^ x2_1_inp);
    assign L3_1 = (Q0_1 ^ x3_1_inp);
    assign b0_preshared_hpc10 = (Q1_0 ^ r1_inp);
    assign b1_preshared_hpc10 = (Q1_1 ^ r1_inp);
    assign p2_hpc10 = (Q0_0_reg & b1_preshared_hpc10_reg);
    assign i1_hpc10 = (p2_hpc10 ^ r2_inp_reg);
    assign p3_hpc10 = (Q0_1_reg & b0_preshared_hpc10_reg);
    assign i2_hpc10 = (p3_hpc10 ^ r2_inp_reg);
    assign p1_hpc10 = (Q0_0_reg & b0_preshared_hpc10_reg);
    assign p4_hpc10 = (Q0_1_reg & b1_preshared_hpc10_reg);
    assign T0_0 = (i1_hpc10_reg ^ p1_hpc10_reg);
    assign T0_1 = (i2_hpc10_reg ^ p4_hpc10_reg);
    assign L10_0 = !L2_0;
    assign L10_1 = !L2_1;
    assign b0_preshared_hpc11 = (Q4_0 ^ r1_inp);
    assign b1_preshared_hpc11 = (Q4_1 ^ r1_inp);
    assign p2_hpc11 = (x1_0_inp_reg & b1_preshared_hpc11_reg);
    assign i1_hpc11 = (p2_hpc11 ^ r2_inp_reg);
    assign p3_hpc11 = (x1_1_inp_reg & b0_preshared_hpc11_reg);
    assign i2_hpc11 = (p3_hpc11 ^ r2_inp_reg);
    assign p1_hpc11 = (x1_0_inp_reg & b0_preshared_hpc11_reg);
    assign p4_hpc11 = (x1_1_inp_reg & b1_preshared_hpc11_reg);
    assign T2_0 = (i1_hpc11_reg ^ p1_hpc11_reg);
    assign T2_1 = (i2_hpc11_reg ^ p4_hpc11_reg);
    assign z329_assgn329 = L2_0;
    assign Q2_0 = (T0_0 ^ z121_assgn121);
    assign L4_0 = (T0_0 ^ T2_0);
    assign z335_assgn335 = L5_0;
    assign Q7_0 = (T0_0 ^ z125_assgn125);
    assign z339_assgn339 = L3_0;
    assign Q6_0 = (L4_0 ^ z127_assgn127);
    assign z343_assgn343 = L2_1;
    assign Q2_1 = (T0_1 ^ z129_assgn129);
    assign L4_1 = (T0_1 ^ T2_1);
    assign z349_assgn349 = L5_1;
    assign Q7_1 = (T0_1 ^ z133_assgn133);
    assign z353_assgn353 = L3_1;
    assign Q6_1 = (L4_1 ^ z135_assgn135);
    assign b0_preshared_hpc12 = (Q3_0 ^ r1_inp);
    assign b1_preshared_hpc12 = (Q3_1 ^ r1_inp);
    assign z361_assgn361 = b1_preshared_hpc12;
    assign p2_hpc12 = (Q2_0 & z141_assgn141);
    assign z365_assgn365 = r2_inp;
    assign i1_hpc12 = (p2_hpc12 ^ z143_assgn143);
    assign z369_assgn369 = b0_preshared_hpc12;
    assign p3_hpc12 = (Q2_1 & z145_assgn145);
    assign z373_assgn373 = r2_inp;
    assign i2_hpc12 = (p3_hpc12 ^ z147_assgn147);
    assign z377_assgn377 = b0_preshared_hpc12;
    assign p1_hpc12 = (Q2_0 & z149_assgn149);
    assign z381_assgn381 = b1_preshared_hpc12;
    assign p4_hpc12 = (Q2_1 & z151_assgn151);
    assign T1_0 = (i1_hpc12_reg ^ p1_hpc12_reg);
    assign T1_1 = (i2_hpc12_reg ^ p4_hpc12_reg);
    assign z389_assgn389 = r1_inp;
    assign b0_preshared_hpc13 = (Q7_0 ^ z157_assgn157);
    assign z393_assgn393 = r1_inp;
    assign b1_preshared_hpc13 = (Q7_1 ^ z159_assgn159);
    assign p2_hpc13 = (Q6_0_reg & b1_preshared_hpc13_reg);
    assign z399_assgn399 = r2_inp;
    assign i1_hpc13 = (p2_hpc13 ^ z163_assgn163);
    assign p3_hpc13 = (Q6_1_reg & b0_preshared_hpc13_reg);
    assign z405_assgn405 = r2_inp;
    assign i2_hpc13 = (p3_hpc13 ^ z167_assgn167);
    assign p1_hpc13 = (Q6_0_reg & b0_preshared_hpc13_reg);
    assign p4_hpc13 = (Q6_1_reg & b1_preshared_hpc13_reg);
    assign T3_0 = (i1_hpc13_reg ^ p1_hpc13_reg);
    assign T3_1 = (i2_hpc13_reg ^ p4_hpc13_reg);
    assign L7_0 = (T0_0_reg ^ T1_0);
    assign z419_assgn419 = L10_0;
    assign L11_0 = (T1_0 ^ z179_assgn179);
    assign L7_1 = (T0_1_reg ^ T1_1);
    assign z425_assgn425 = L10_1;
    assign L11_1 = (T1_1 ^ z183_assgn183);
    assign Y0_01 = (L7_0 ^ T2_0_reg);
    assign z431_assgn431 = L8_0;
    assign Y1_01 = (z188_assgn188 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1_reg);
    assign z437_assgn437 = L8_1;
    assign Y1_11 = (z192_assgn192 ^ T3_1);
    assign z441_assgn441 = x3_0_inp;
    assign z1_assgn1 = (z194_assgn194 ^ Y0_01);
    assign z445_assgn445 = z1_assgn1;
    assign z3_assgn3 = (L7_0_reg ^ Y1_01);
    assign z5_assgn5 = (L11_0 ^ T2_0_reg);
    assign z453_assgn453 = z5_assgn5;
    assign z455_assgn455 = L5_0;
    assign z7_assgn7 = (T2_0 ^ z205_assgn205);
    assign z459_assgn459 = z7_assgn7;
    assign z461_assgn461 = x3_1_inp;
    assign z9_assgn9 = (z210_assgn210 ^ Y0_11);
    assign z465_assgn465 = z9_assgn9;
    assign z11_assgn11 = (L7_1_reg ^ Y1_11);
    assign z13_assgn13 = (L11_1 ^ T2_1_reg);
    assign z473_assgn473 = z13_assgn13;
    assign z475_assgn475 = L5_1;
    assign z15_assgn15 = (T2_1 ^ z221_assgn221);
    assign z479_assgn479 = z15_assgn15;

    always @(posedge clk) begin
        Q0_0_reg <= Q0_0;
        b1_preshared_hpc10_reg <= b1_preshared_hpc10;
        r2_inp_reg <= r2_inp;
        Q0_1_reg <= Q0_1;
        b0_preshared_hpc10_reg <= b0_preshared_hpc10;
        i1_hpc10_reg <= i1_hpc10;
        p1_hpc10_reg <= p1_hpc10;
        i2_hpc10_reg <= i2_hpc10;
        p4_hpc10_reg <= p4_hpc10;
        x1_0_inp_reg <= x1_0_inp;
        b1_preshared_hpc11_reg <= b1_preshared_hpc11;
        x1_1_inp_reg <= x1_1_inp;
        b0_preshared_hpc11_reg <= b0_preshared_hpc11;
        i1_hpc11_reg <= i1_hpc11;
        p1_hpc11_reg <= p1_hpc11;
        i2_hpc11_reg <= i2_hpc11;
        p4_hpc11_reg <= p4_hpc11;
        z329_assgn3290 <= z329_assgn329;
        z121_assgn121 <= z329_assgn3290;
        z335_assgn3350 <= z335_assgn335;
        z125_assgn125 <= z335_assgn3350;
        z339_assgn3390 <= z339_assgn339;
        z127_assgn127 <= z339_assgn3390;
        z343_assgn3430 <= z343_assgn343;
        z129_assgn129 <= z343_assgn3430;
        z349_assgn3490 <= z349_assgn349;
        z133_assgn133 <= z349_assgn3490;
        z353_assgn3530 <= z353_assgn353;
        z135_assgn135 <= z353_assgn3530;
        z361_assgn3610 <= z361_assgn361;
        z141_assgn141 <= z361_assgn3610;
        z365_assgn3650 <= z365_assgn365;
        z143_assgn143 <= z365_assgn3650;
        z369_assgn3690 <= z369_assgn369;
        z145_assgn145 <= z369_assgn3690;
        z373_assgn3730 <= z373_assgn373;
        z147_assgn147 <= z373_assgn3730;
        z377_assgn3770 <= z377_assgn377;
        z149_assgn149 <= z377_assgn3770;
        z381_assgn3810 <= z381_assgn381;
        z151_assgn151 <= z381_assgn3810;
        i1_hpc12_reg <= i1_hpc12;
        p1_hpc12_reg <= p1_hpc12;
        i2_hpc12_reg <= i2_hpc12;
        p4_hpc12_reg <= p4_hpc12;
        z389_assgn3890 <= z389_assgn389;
        z157_assgn157 <= z389_assgn3890;
        z393_assgn3930 <= z393_assgn393;
        z159_assgn159 <= z393_assgn3930;
        Q6_0_reg <= Q6_0;
        b1_preshared_hpc13_reg <= b1_preshared_hpc13;
        z399_assgn3990 <= z399_assgn399;
        z399_assgn3991 <= z399_assgn3990;
        z163_assgn163 <= z399_assgn3991;
        Q6_1_reg <= Q6_1;
        b0_preshared_hpc13_reg <= b0_preshared_hpc13;
        z405_assgn4050 <= z405_assgn405;
        z405_assgn4051 <= z405_assgn4050;
        z167_assgn167 <= z405_assgn4051;
        i1_hpc13_reg <= i1_hpc13;
        p1_hpc13_reg <= p1_hpc13;
        i2_hpc13_reg <= i2_hpc13;
        p4_hpc13_reg <= p4_hpc13;
        T0_0_reg <= T0_0;
        z419_assgn4190 <= z419_assgn419;
        z419_assgn4191 <= z419_assgn4190;
        z179_assgn179 <= z419_assgn4191;
        T0_1_reg <= T0_1;
        z425_assgn4250 <= z425_assgn425;
        z425_assgn4251 <= z425_assgn4250;
        z183_assgn183 <= z425_assgn4251;
        T2_0_reg <= T2_0;
        z431_assgn4310 <= z431_assgn431;
        z431_assgn4311 <= z431_assgn4310;
        z431_assgn4312 <= z431_assgn4311;
        z188_assgn188 <= z431_assgn4312;
        T2_1_reg <= T2_1;
        z437_assgn4370 <= z437_assgn437;
        z437_assgn4371 <= z437_assgn4370;
        z437_assgn4372 <= z437_assgn4371;
        z192_assgn192 <= z437_assgn4372;
        z441_assgn4410 <= z441_assgn441;
        z441_assgn4411 <= z441_assgn4410;
        z194_assgn194 <= z441_assgn4411;
        z445_assgn4450 <= z445_assgn445;
        Y0_0 <= z445_assgn4450;
        L7_0_reg <= L7_0;
        Y1_0 <= z3_assgn3;
        z453_assgn4530 <= z453_assgn453;
        Y2_0 <= z453_assgn4530;
        z455_assgn4550 <= z455_assgn455;
        z205_assgn205 <= z455_assgn4550;
        z459_assgn4590 <= z459_assgn459;
        z459_assgn4591 <= z459_assgn4590;
        Y3_0 <= z459_assgn4591;
        z461_assgn4610 <= z461_assgn461;
        z461_assgn4611 <= z461_assgn4610;
        z210_assgn210 <= z461_assgn4611;
        z465_assgn4650 <= z465_assgn465;
        Y0_1 <= z465_assgn4650;
        L7_1_reg <= L7_1;
        Y1_1 <= z11_assgn11;
        z473_assgn4730 <= z473_assgn473;
        Y2_1 <= z473_assgn4730;
        z475_assgn4750 <= z475_assgn475;
        z221_assgn221 <= z475_assgn4750;
        z479_assgn4790 <= z479_assgn479;
        z479_assgn4791 <= z479_assgn4790;
        Y3_1 <= z479_assgn4791;
    end

endmodule

