module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    wire x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    wire x3_1_inp;
    wire r_inp;
    wire L0_0;
    wire L1_0;
    wire L8_0;
    wire L5_0;
    wire L0_1;
    wire L1_1;
    wire L8_1;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire L2_0;
    wire L3_0;
    wire L2_1;
    wire L3_1;
    wire a0_neg_hpc20;
    wire a1_neg_hpc20;
    reg a0_neg_hpc20_reg;
    reg r_inp_reg;
    wire u0_hpc20;
    reg a1_neg_hpc20_reg;
    wire u1_hpc20;
    wire v0_hpc20;
    wire v1_hpc20;
    reg Q0_0_reg;
    reg Q1_0_reg;
    wire p0_hpc20;
    reg v1_hpc20_reg;
    wire p1_hpc20;
    reg u0_hpc20_reg;
    reg p1_hpc20_reg;
    wire p01_hpc20;
    reg p0_hpc20_reg;
    wire T0_0;
    reg Q0_1_reg;
    reg Q1_1_reg;
    wire p2_hpc20;
    reg v0_hpc20_reg;
    wire p3_hpc20;
    reg u1_hpc20_reg;
    reg p3_hpc20_reg;
    wire p23_hpc20;
    reg p2_hpc20_reg;
    wire T0_1;
    wire L10_0;
    wire L10_1;
    wire a0_neg_hpc21;
    wire a1_neg_hpc21;
    reg a0_neg_hpc21_reg;
    wire u0_hpc21;
    reg a1_neg_hpc21_reg;
    wire u1_hpc21;
    wire v0_hpc21;
    wire v1_hpc21;
    reg x1_0_inp_reg;
    reg Q4_0_reg;
    wire p0_hpc21;
    reg v1_hpc21_reg;
    wire p1_hpc21;
    reg u0_hpc21_reg;
    reg p1_hpc21_reg;
    wire p01_hpc21;
    reg p0_hpc21_reg;
    wire T2_0;
    reg x1_1_inp_reg;
    reg Q4_1_reg;
    wire p2_hpc21;
    reg v0_hpc21_reg;
    wire p3_hpc21;
    reg u1_hpc21_reg;
    reg p3_hpc21_reg;
    wire p23_hpc21;
    reg p2_hpc21_reg;
    wire T2_1;
    wire z373_assgn373;
    reg z373_assgn3730;
    reg z135_assgn135;
    wire Q2_0;
    wire L4_0;
    wire z379_assgn379;
    reg z379_assgn3790;
    reg z139_assgn139;
    wire Q7_0;
    wire z383_assgn383;
    reg z383_assgn3830;
    reg z141_assgn141;
    wire Q6_0;
    wire z387_assgn387;
    reg z387_assgn3870;
    reg z143_assgn143;
    wire Q2_1;
    wire L4_1;
    wire z393_assgn393;
    reg z393_assgn3930;
    reg z147_assgn147;
    wire Q7_1;
    wire z397_assgn397;
    reg z397_assgn3970;
    reg z149_assgn149;
    wire Q6_1;
    wire a0_neg_hpc22;
    wire a1_neg_hpc22;
    wire z405_assgn405;
    reg z405_assgn4050;
    reg z155_assgn155;
    wire u0_hpc22;
    wire z409_assgn409;
    reg z409_assgn4090;
    reg z157_assgn157;
    wire u1_hpc22;
    wire v0_hpc22;
    wire v1_hpc22;
    wire z417_assgn417;
    reg z417_assgn4170;
    reg z163_assgn163;
    wire p0_hpc22;
    wire z421_assgn421;
    reg z421_assgn4210;
    reg z165_assgn165;
    wire p1_hpc22;
    reg u0_hpc22_reg;
    reg p1_hpc22_reg;
    wire p01_hpc22;
    reg p0_hpc22_reg;
    wire T1_0;
    wire z429_assgn429;
    reg z429_assgn4290;
    reg z171_assgn171;
    wire p2_hpc22;
    wire z433_assgn433;
    reg z433_assgn4330;
    reg z173_assgn173;
    wire p3_hpc22;
    reg u1_hpc22_reg;
    reg p3_hpc22_reg;
    wire p23_hpc22;
    reg p2_hpc22_reg;
    wire T1_1;
    wire a0_neg_hpc23;
    wire a1_neg_hpc23;
    wire z445_assgn445;
    reg z445_assgn4450;
    reg z183_assgn183;
    wire u0_hpc23;
    wire z449_assgn449;
    reg z449_assgn4490;
    reg z185_assgn185;
    wire u1_hpc23;
    wire z453_assgn453;
    reg z453_assgn4530;
    reg z187_assgn187;
    wire v0_hpc23;
    wire z457_assgn457;
    reg z457_assgn4570;
    reg z189_assgn189;
    wire v1_hpc23;
    reg Q6_0_reg;
    reg Q7_0_reg;
    wire p0_hpc23;
    reg v1_hpc23_reg;
    wire p1_hpc23;
    wire z465_assgn465;
    reg z465_assgn4650;
    reg z196_assgn196;
    reg p1_hpc23_reg;
    wire p01_hpc23;
    reg p0_hpc23_reg;
    wire T3_0;
    reg Q6_1_reg;
    reg Q7_1_reg;
    wire p2_hpc23;
    reg v0_hpc23_reg;
    wire p3_hpc23;
    wire z475_assgn475;
    reg z475_assgn4750;
    reg z204_assgn204;
    reg p3_hpc23_reg;
    wire p23_hpc23;
    reg p2_hpc23_reg;
    wire T3_1;
    reg T0_0_reg;
    wire L7_0;
    wire z483_assgn483;
    reg z483_assgn4830;
    reg z483_assgn4831;
    reg z209_assgn209;
    wire L11_0;
    reg T0_1_reg;
    wire L7_1;
    wire z489_assgn489;
    reg z489_assgn4890;
    reg z489_assgn4891;
    reg z213_assgn213;
    wire L11_1;
    reg T2_0_reg;
    wire Y0_01;
    wire z495_assgn495;
    reg z495_assgn4950;
    reg z495_assgn4951;
    reg z495_assgn4952;
    reg z218_assgn218;
    wire Y1_01;
    reg T2_1_reg;
    wire Y0_11;
    wire z501_assgn501;
    reg z501_assgn5010;
    reg z501_assgn5011;
    reg z501_assgn5012;
    reg z222_assgn222;
    wire Y1_11;
    wire z505_assgn505;
    reg z505_assgn5050;
    reg z505_assgn5051;
    reg z224_assgn224;
    wire z1_assgn1;
    wire z509_assgn509;
    reg z509_assgn5090;
    reg L7_0_reg;
    wire z3_assgn3;
    wire z5_assgn5;
    wire z517_assgn517;
    reg z517_assgn5170;
    wire z519_assgn519;
    reg z519_assgn5190;
    reg z235_assgn235;
    wire z7_assgn7;
    wire z523_assgn523;
    reg z523_assgn5230;
    reg z523_assgn5231;
    wire z525_assgn525;
    reg z525_assgn5250;
    reg z525_assgn5251;
    reg z240_assgn240;
    wire z9_assgn9;
    wire z529_assgn529;
    reg z529_assgn5290;
    reg L7_1_reg;
    wire z11_assgn11;
    wire z13_assgn13;
    wire z537_assgn537;
    reg z537_assgn5370;
    wire z539_assgn539;
    reg z539_assgn5390;
    reg z251_assgn251;
    wire z15_assgn15;
    wire z543_assgn543;
    reg z543_assgn5430;
    reg z543_assgn5431;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign x3_0_inp = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign x3_1_inp = x3_1;
    assign r_inp = r;
    assign L0_0 = (x1_0_inp ^ x2_0_inp);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign L8_0 = (x2_0_inp ^ x0_0_inp);
    assign L5_0 = (x0_0_inp ^ x3_0_inp);
    assign L0_1 = (x1_1_inp ^ x2_1_inp);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign L8_1 = (x2_1_inp ^ x0_1_inp);
    assign L5_1 = (x0_1_inp ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !x2_0_inp;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !x2_1_inp;
    assign L2_0 = (Q1_0 ^ x2_0_inp);
    assign L3_0 = (Q0_0 ^ x3_0_inp);
    assign L2_1 = (Q1_1 ^ x2_1_inp);
    assign L3_1 = (Q0_1 ^ x3_1_inp);
    assign a0_neg_hpc20 = !Q0_0;
    assign a1_neg_hpc20 = !Q0_1;
    assign u0_hpc20 = (a0_neg_hpc20_reg & r_inp_reg);
    assign u1_hpc20 = (a1_neg_hpc20_reg & r_inp_reg);
    assign v0_hpc20 = (Q1_0 ^ r_inp);
    assign v1_hpc20 = (Q1_1 ^ r_inp);
    assign p0_hpc20 = (Q0_0_reg & Q1_0_reg);
    assign p1_hpc20 = (Q0_0_reg & v1_hpc20_reg);
    assign p01_hpc20 = (u0_hpc20_reg ^ p1_hpc20_reg);
    assign T0_0 = (p0_hpc20_reg ^ p01_hpc20);
    assign p2_hpc20 = (Q0_1_reg & Q1_1_reg);
    assign p3_hpc20 = (Q0_1_reg & v0_hpc20_reg);
    assign p23_hpc20 = (u1_hpc20_reg ^ p3_hpc20_reg);
    assign T0_1 = (p2_hpc20_reg ^ p23_hpc20);
    assign L10_0 = !L2_0;
    assign L10_1 = !L2_1;
    assign a0_neg_hpc21 = !x1_0_inp;
    assign a1_neg_hpc21 = !x1_1_inp;
    assign u0_hpc21 = (a0_neg_hpc21_reg & r_inp_reg);
    assign u1_hpc21 = (a1_neg_hpc21_reg & r_inp_reg);
    assign v0_hpc21 = (Q4_0 ^ r_inp);
    assign v1_hpc21 = (Q4_1 ^ r_inp);
    assign p0_hpc21 = (x1_0_inp_reg & Q4_0_reg);
    assign p1_hpc21 = (x1_0_inp_reg & v1_hpc21_reg);
    assign p01_hpc21 = (u0_hpc21_reg ^ p1_hpc21_reg);
    assign T2_0 = (p0_hpc21_reg ^ p01_hpc21);
    assign p2_hpc21 = (x1_1_inp_reg & Q4_1_reg);
    assign p3_hpc21 = (x1_1_inp_reg & v0_hpc21_reg);
    assign p23_hpc21 = (u1_hpc21_reg ^ p3_hpc21_reg);
    assign T2_1 = (p2_hpc21_reg ^ p23_hpc21);
    assign z373_assgn373 = L2_0;
    assign Q2_0 = (T0_0 ^ z135_assgn135);
    assign L4_0 = (T0_0 ^ T2_0);
    assign z379_assgn379 = L5_0;
    assign Q7_0 = (T0_0 ^ z139_assgn139);
    assign z383_assgn383 = L3_0;
    assign Q6_0 = (L4_0 ^ z141_assgn141);
    assign z387_assgn387 = L2_1;
    assign Q2_1 = (T0_1 ^ z143_assgn143);
    assign L4_1 = (T0_1 ^ T2_1);
    assign z393_assgn393 = L5_1;
    assign Q7_1 = (T0_1 ^ z147_assgn147);
    assign z397_assgn397 = L3_1;
    assign Q6_1 = (L4_1 ^ z149_assgn149);
    assign a0_neg_hpc22 = !Q2_0;
    assign a1_neg_hpc22 = !Q2_1;
    assign z405_assgn405 = r_inp;
    assign u0_hpc22 = (a0_neg_hpc22 & z155_assgn155);
    assign z409_assgn409 = r_inp;
    assign u1_hpc22 = (a1_neg_hpc22 & z157_assgn157);
    assign v0_hpc22 = (Q3_0 ^ r_inp);
    assign v1_hpc22 = (Q3_1 ^ r_inp);
    assign z417_assgn417 = Q3_0;
    assign p0_hpc22 = (Q2_0 & z163_assgn163);
    assign z421_assgn421 = v1_hpc22;
    assign p1_hpc22 = (Q2_0 & z165_assgn165);
    assign p01_hpc22 = (u0_hpc22_reg ^ p1_hpc22_reg);
    assign T1_0 = (p0_hpc22_reg ^ p01_hpc22);
    assign z429_assgn429 = Q3_1;
    assign p2_hpc22 = (Q2_1 & z171_assgn171);
    assign z433_assgn433 = v0_hpc22;
    assign p3_hpc22 = (Q2_1 & z173_assgn173);
    assign p23_hpc22 = (u1_hpc22_reg ^ p3_hpc22_reg);
    assign T1_1 = (p2_hpc22_reg ^ p23_hpc22);
    assign a0_neg_hpc23 = !Q6_0;
    assign a1_neg_hpc23 = !Q6_1;
    assign z445_assgn445 = r_inp;
    assign u0_hpc23 = (a0_neg_hpc23 & z183_assgn183);
    assign z449_assgn449 = r_inp;
    assign u1_hpc23 = (a1_neg_hpc23 & z185_assgn185);
    assign z453_assgn453 = r_inp;
    assign v0_hpc23 = (Q7_0 ^ z187_assgn187);
    assign z457_assgn457 = r_inp;
    assign v1_hpc23 = (Q7_1 ^ z189_assgn189);
    assign p0_hpc23 = (Q6_0_reg & Q7_0_reg);
    assign p1_hpc23 = (Q6_0_reg & v1_hpc23_reg);
    assign z465_assgn465 = u0_hpc23;
    assign p01_hpc23 = (z196_assgn196 ^ p1_hpc23_reg);
    assign T3_0 = (p0_hpc23_reg ^ p01_hpc23);
    assign p2_hpc23 = (Q6_1_reg & Q7_1_reg);
    assign p3_hpc23 = (Q6_1_reg & v0_hpc23_reg);
    assign z475_assgn475 = u1_hpc23;
    assign p23_hpc23 = (z204_assgn204 ^ p3_hpc23_reg);
    assign T3_1 = (p2_hpc23_reg ^ p23_hpc23);
    assign L7_0 = (T0_0_reg ^ T1_0);
    assign z483_assgn483 = L10_0;
    assign L11_0 = (T1_0 ^ z209_assgn209);
    assign L7_1 = (T0_1_reg ^ T1_1);
    assign z489_assgn489 = L10_1;
    assign L11_1 = (T1_1 ^ z213_assgn213);
    assign Y0_01 = (L7_0 ^ T2_0_reg);
    assign z495_assgn495 = L8_0;
    assign Y1_01 = (z218_assgn218 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1_reg);
    assign z501_assgn501 = L8_1;
    assign Y1_11 = (z222_assgn222 ^ T3_1);
    assign z505_assgn505 = x3_0_inp;
    assign z1_assgn1 = (z224_assgn224 ^ Y0_01);
    assign z509_assgn509 = z1_assgn1;
    assign z3_assgn3 = (L7_0_reg ^ Y1_01);
    assign z5_assgn5 = (L11_0 ^ T2_0_reg);
    assign z517_assgn517 = z5_assgn5;
    assign z519_assgn519 = L5_0;
    assign z7_assgn7 = (T2_0 ^ z235_assgn235);
    assign z523_assgn523 = z7_assgn7;
    assign z525_assgn525 = x3_1_inp;
    assign z9_assgn9 = (z240_assgn240 ^ Y0_11);
    assign z529_assgn529 = z9_assgn9;
    assign z11_assgn11 = (L7_1_reg ^ Y1_11);
    assign z13_assgn13 = (L11_1 ^ T2_1_reg);
    assign z537_assgn537 = z13_assgn13;
    assign z539_assgn539 = L5_1;
    assign z15_assgn15 = (T2_1 ^ z251_assgn251);
    assign z543_assgn543 = z15_assgn15;

    always @(posedge clk) begin
        a0_neg_hpc20_reg <= a0_neg_hpc20;
        r_inp_reg <= r_inp;
        a1_neg_hpc20_reg <= a1_neg_hpc20;
        Q0_0_reg <= Q0_0;
        Q1_0_reg <= Q1_0;
        v1_hpc20_reg <= v1_hpc20;
        u0_hpc20_reg <= u0_hpc20;
        p1_hpc20_reg <= p1_hpc20;
        p0_hpc20_reg <= p0_hpc20;
        Q0_1_reg <= Q0_1;
        Q1_1_reg <= Q1_1;
        v0_hpc20_reg <= v0_hpc20;
        u1_hpc20_reg <= u1_hpc20;
        p3_hpc20_reg <= p3_hpc20;
        p2_hpc20_reg <= p2_hpc20;
        a0_neg_hpc21_reg <= a0_neg_hpc21;
        a1_neg_hpc21_reg <= a1_neg_hpc21;
        x1_0_inp_reg <= x1_0_inp;
        Q4_0_reg <= Q4_0;
        v1_hpc21_reg <= v1_hpc21;
        u0_hpc21_reg <= u0_hpc21;
        p1_hpc21_reg <= p1_hpc21;
        p0_hpc21_reg <= p0_hpc21;
        x1_1_inp_reg <= x1_1_inp;
        Q4_1_reg <= Q4_1;
        v0_hpc21_reg <= v0_hpc21;
        u1_hpc21_reg <= u1_hpc21;
        p3_hpc21_reg <= p3_hpc21;
        p2_hpc21_reg <= p2_hpc21;
        z373_assgn3730 <= z373_assgn373;
        z135_assgn135 <= z373_assgn3730;
        z379_assgn3790 <= z379_assgn379;
        z139_assgn139 <= z379_assgn3790;
        z383_assgn3830 <= z383_assgn383;
        z141_assgn141 <= z383_assgn3830;
        z387_assgn3870 <= z387_assgn387;
        z143_assgn143 <= z387_assgn3870;
        z393_assgn3930 <= z393_assgn393;
        z147_assgn147 <= z393_assgn3930;
        z397_assgn3970 <= z397_assgn397;
        z149_assgn149 <= z397_assgn3970;
        z405_assgn4050 <= z405_assgn405;
        z155_assgn155 <= z405_assgn4050;
        z409_assgn4090 <= z409_assgn409;
        z157_assgn157 <= z409_assgn4090;
        z417_assgn4170 <= z417_assgn417;
        z163_assgn163 <= z417_assgn4170;
        z421_assgn4210 <= z421_assgn421;
        z165_assgn165 <= z421_assgn4210;
        u0_hpc22_reg <= u0_hpc22;
        p1_hpc22_reg <= p1_hpc22;
        p0_hpc22_reg <= p0_hpc22;
        z429_assgn4290 <= z429_assgn429;
        z171_assgn171 <= z429_assgn4290;
        z433_assgn4330 <= z433_assgn433;
        z173_assgn173 <= z433_assgn4330;
        u1_hpc22_reg <= u1_hpc22;
        p3_hpc22_reg <= p3_hpc22;
        p2_hpc22_reg <= p2_hpc22;
        z445_assgn4450 <= z445_assgn445;
        z183_assgn183 <= z445_assgn4450;
        z449_assgn4490 <= z449_assgn449;
        z185_assgn185 <= z449_assgn4490;
        z453_assgn4530 <= z453_assgn453;
        z187_assgn187 <= z453_assgn4530;
        z457_assgn4570 <= z457_assgn457;
        z189_assgn189 <= z457_assgn4570;
        Q6_0_reg <= Q6_0;
        Q7_0_reg <= Q7_0;
        v1_hpc23_reg <= v1_hpc23;
        z465_assgn4650 <= z465_assgn465;
        z196_assgn196 <= z465_assgn4650;
        p1_hpc23_reg <= p1_hpc23;
        p0_hpc23_reg <= p0_hpc23;
        Q6_1_reg <= Q6_1;
        Q7_1_reg <= Q7_1;
        v0_hpc23_reg <= v0_hpc23;
        z475_assgn4750 <= z475_assgn475;
        z204_assgn204 <= z475_assgn4750;
        p3_hpc23_reg <= p3_hpc23;
        p2_hpc23_reg <= p2_hpc23;
        T0_0_reg <= T0_0;
        z483_assgn4830 <= z483_assgn483;
        z483_assgn4831 <= z483_assgn4830;
        z209_assgn209 <= z483_assgn4831;
        T0_1_reg <= T0_1;
        z489_assgn4890 <= z489_assgn489;
        z489_assgn4891 <= z489_assgn4890;
        z213_assgn213 <= z489_assgn4891;
        T2_0_reg <= T2_0;
        z495_assgn4950 <= z495_assgn495;
        z495_assgn4951 <= z495_assgn4950;
        z495_assgn4952 <= z495_assgn4951;
        z218_assgn218 <= z495_assgn4952;
        T2_1_reg <= T2_1;
        z501_assgn5010 <= z501_assgn501;
        z501_assgn5011 <= z501_assgn5010;
        z501_assgn5012 <= z501_assgn5011;
        z222_assgn222 <= z501_assgn5012;
        z505_assgn5050 <= z505_assgn505;
        z505_assgn5051 <= z505_assgn5050;
        z224_assgn224 <= z505_assgn5051;
        z509_assgn5090 <= z509_assgn509;
        Y0_0 <= z509_assgn5090;
        L7_0_reg <= L7_0;
        Y1_0 <= z3_assgn3;
        z517_assgn5170 <= z517_assgn517;
        Y2_0 <= z517_assgn5170;
        z519_assgn5190 <= z519_assgn519;
        z235_assgn235 <= z519_assgn5190;
        z523_assgn5230 <= z523_assgn523;
        z523_assgn5231 <= z523_assgn5230;
        Y3_0 <= z523_assgn5231;
        z525_assgn5250 <= z525_assgn525;
        z525_assgn5251 <= z525_assgn5250;
        z240_assgn240 <= z525_assgn5251;
        z529_assgn5290 <= z529_assgn529;
        Y0_1 <= z529_assgn5290;
        L7_1_reg <= L7_1;
        Y1_1 <= z11_assgn11;
        z537_assgn5370 <= z537_assgn537;
        Y2_1 <= z537_assgn5370;
        z539_assgn5390 <= z539_assgn539;
        z251_assgn251 <= z539_assgn5390;
        z543_assgn5430 <= z543_assgn543;
        z543_assgn5431 <= z543_assgn5430;
        Y3_1 <= z543_assgn5431;
    end

endmodule

