module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    r6,
    r7,
    r8,
    r9,
    r10,
    r11,
    r12,
    r13,
    r14,
    r15,
    r16,
    r17,
    r18,
    r19,
    r20,
    r21,
    r22,
    r23,
    r24,
    r25,
    r26,
    r27,
    r28,
    r29,
    r30,
    r31,
    r32,
    r33,
    r34,
    r35,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1
);
//INPUTS
    input clk;
    input [7:0]  t0;
    input [7:0]  t1;
    input [7:0]  r0;
    input [7:0]  r1;
    input [7:0]  r2;
    input [7:0]  r3;
    input [7:0]  r4;
    input [7:0]  r5;
    input [7:0]  r6;
    input [7:0]  r7;
    input [7:0]  r8;
    input [7:0]  r9;
    input [7:0]  r10;
    input [7:0]  r11;
    input [7:0]  r12;
    input [7:0]  r13;
    input [7:0]  r14;
    input [7:0]  r15;
    input [7:0]  r16;
    input [7:0]  r17;
    input [7:0]  r18;
    input [7:0]  r19;
    input [7:0]  r20;
    input [7:0]  r21;
    input [7:0]  r22;
    input [7:0]  r23;
    input [7:0]  r24;
    input [7:0]  r25;
    input [7:0]  r26;
    input [7:0]  r27;
    input [7:0]  r28;
    input [7:0]  r29;
    input [7:0]  r30;
    input [7:0]  r31;
    input [7:0]  r32;
    input [7:0]  r33;
    input [7:0]  r34;
    input [7:0]  r35;
    input [7:0]  dec_0;
    input [7:0]  dec_1;
    input [7:0]  dec_255;
    input [7:0]  dec_169;
    input [7:0]  dec_129;
    input [7:0]  dec_9;
    input [7:0]  dec_72;
    input [7:0]  dec_242;
    input [7:0]  dec_243;
    input [7:0]  dec_152;
    input [7:0]  dec_240;
    input [7:0]  dec_4;
    input [7:0]  dec_15;
    input [7:0]  dec_12;
    input [7:0]  dec_2;
    input [7:0]  dec_3;
    input [7:0]  dec_16;
    input [7:0]  dec_36;
    input [7:0]  dec_220;
    input [7:0]  dec_11;
    input [7:0]  dec_158;
    input [7:0]  dec_45;
    input [7:0]  dec_88;
    input [7:0]  dec_99;
//OUTPUTS
    output reg [7:0]  y0;
    output reg [7:0]  y1;
//Intermediate values
    wire [7:0] dec_99_inp;
    wire [7:0] dec_88_inp;
    wire [7:0] dec_45_inp;
    wire [7:0] dec_158_inp;
    wire [7:0] dec_11_inp;
    wire [7:0] dec_220_inp;
    wire [7:0] dec_36_inp;
    wire [7:0] dec_16_inp;
    wire [7:0] dec_3_inp;
    wire [7:0] dec_2_inp;
    wire [7:0] dec_12_inp;
    wire [7:0] dec_15_inp;
    wire [7:0] dec_4_inp;
    wire [7:0] dec_240_inp;
    wire [7:0] dec_152_inp;
    wire [7:0] dec_243_inp;
    wire [7:0] dec_242_inp;
    wire [7:0] dec_72_inp;
    wire [7:0] dec_9_inp;
    wire [7:0] dec_129_inp;
    wire [7:0] dec_169_inp;
    wire [7:0] dec_255_inp;
    wire [7:0] dec_1_inp;
    wire [7:0] dec_0_inp;
    wire [7:0] t0_inp;
    wire [7:0] t1_inp;
    wire [7:0] r0_inp;
    wire [7:0] r1_inp;
    wire [7:0] r2_inp;
    wire [7:0] r3_inp;
    wire [7:0] r4_inp;
    wire [7:0] r5_inp;
    wire [7:0] r6_inp;
    wire [7:0] r7_inp;
    wire [7:0] r8_inp;
    wire [7:0] r9_inp;
    wire [7:0] r10_inp;
    wire [7:0] r11_inp;
    wire [7:0] r12_inp;
    wire [7:0] r13_inp;
    wire [7:0] r14_inp;
    wire [7:0] r15_inp;
    wire [7:0] r16_inp;
    wire [7:0] r17_inp;
    wire [7:0] r18_inp;
    wire [7:0] r19_inp;
    wire [7:0] r20_inp;
    wire [7:0] r21_inp;
    wire [7:0] r22_inp;
    wire [7:0] r23_inp;
    wire [7:0] r24_inp;
    wire [7:0] r25_inp;
    wire [7:0] r26_inp;
    wire [7:0] r27_inp;
    wire [7:0] r28_inp;
    wire [7:0] r29_inp;
    wire [7:0] r30_inp;
    wire [7:0] r31_inp;
    wire [7:0] r32_inp;
    wire [7:0] r33_inp;
    wire [7:0] r34_inp;
    wire [7:0] r35_inp;
    wire [7:0] y_G256_newbasis0;
    wire [7:0] tempy1_G256_newbasis0;
    wire [7:0] cond1_G256_newbasis0;
    wire [7:0] negCond1_G256_newbasis0;
    wire [7:0] yxorb1_G256_newbasis0;
    wire [7:0] ny1_G256_newbasis0;
    wire [7:0] tempyIntoNegCond1_G256_newbasis0;
    wire [7:0] y1_G256_newbasis0;
    wire [7:0] x1_G256_newbasis0;
    wire [7:0] tempy2_G256_newbasis0;
    wire [7:0] cond2_G256_newbasis0;
    wire [7:0] negCond2_G256_newbasis0;
    wire [7:0] yxorb2_G256_newbasis0;
    wire [7:0] ny2_G256_newbasis0;
    wire [7:0] tempyIntoNegCond2_G256_newbasis0;
    wire [7:0] y2_G256_newbasis0;
    wire [7:0] x2_G256_newbasis0;
    wire [7:0] tempy3_G256_newbasis0;
    wire [7:0] cond3_G256_newbasis0;
    wire [7:0] negCond3_G256_newbasis0;
    wire [7:0] yxorb3_G256_newbasis0;
    wire [7:0] ny3_G256_newbasis0;
    wire [7:0] tempyIntoNegCond3_G256_newbasis0;
    wire [7:0] y3_G256_newbasis0;
    wire [7:0] x3_G256_newbasis0;
    wire [7:0] tempy4_G256_newbasis0;
    wire [7:0] cond4_G256_newbasis0;
    wire [7:0] negCond4_G256_newbasis0;
    wire [7:0] yxorb4_G256_newbasis0;
    wire [7:0] ny4_G256_newbasis0;
    wire [7:0] tempyIntoNegCond4_G256_newbasis0;
    wire [7:0] y4_G256_newbasis0;
    wire [7:0] x4_G256_newbasis0;
    wire [7:0] tempy5_G256_newbasis0;
    wire [7:0] cond5_G256_newbasis0;
    wire [7:0] negCond5_G256_newbasis0;
    wire [7:0] yxorb5_G256_newbasis0;
    wire [7:0] ny5_G256_newbasis0;
    wire [7:0] tempyIntoNegCond5_G256_newbasis0;
    wire [7:0] y5_G256_newbasis0;
    wire [7:0] x5_G256_newbasis0;
    wire [7:0] tempy6_G256_newbasis0;
    wire [7:0] cond6_G256_newbasis0;
    wire [7:0] negCond6_G256_newbasis0;
    wire [7:0] yxorb6_G256_newbasis0;
    wire [7:0] ny6_G256_newbasis0;
    wire [7:0] tempyIntoNegCond6_G256_newbasis0;
    wire [7:0] y6_G256_newbasis0;
    wire [7:0] x6_G256_newbasis0;
    wire [7:0] tempy7_G256_newbasis0;
    wire [7:0] cond7_G256_newbasis0;
    wire [7:0] negCond7_G256_newbasis0;
    wire [7:0] yxorb7_G256_newbasis0;
    wire [7:0] ny7_G256_newbasis0;
    wire [7:0] tempyIntoNegCond7_G256_newbasis0;
    wire [7:0] y7_G256_newbasis0;
    wire [7:0] x7_G256_newbasis0;
    wire [7:0] tempy8_G256_newbasis0;
    wire [7:0] cond8_G256_newbasis0;
    wire [7:0] negCond8_G256_newbasis0;
    wire [7:0] yxorb8_G256_newbasis0;
    wire [7:0] ny8_G256_newbasis0;
    wire [7:0] tempyIntoNegCond8_G256_newbasis0;
    wire [7:0] y8_G256_newbasis0;
    wire [7:0] z3153_assgn3153;
    reg [7:0] z3153_assgn31530;
    reg [7:0] z3153_assgn31531;
    reg [7:0] z3153_assgn31532;
    reg [7:0] z3153_assgn31533;
    reg [7:0] z3153_assgn31534;
    reg [7:0] x8_G256_newbasis0;
    wire [7:0] t2;
    wire [7:0] z_y_G256_newbasis0;
    wire [7:0] z_tempy1_G256_newbasis0;
    wire [7:0] z_cond1_G256_newbasis0;
    wire [7:0] z_negCond1_G256_newbasis0;
    wire [7:0] z_yxorb1_G256_newbasis0;
    wire [7:0] z_ny1_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond1_G256_newbasis0;
    wire [7:0] z_y1_G256_newbasis0;
    wire [7:0] z_x1_G256_newbasis0;
    wire [7:0] z_tempy2_G256_newbasis0;
    wire [7:0] z_cond2_G256_newbasis0;
    wire [7:0] z_negCond2_G256_newbasis0;
    wire [7:0] z_yxorb2_G256_newbasis0;
    wire [7:0] z_ny2_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond2_G256_newbasis0;
    wire [7:0] z_y2_G256_newbasis0;
    wire [7:0] z_x2_G256_newbasis0;
    wire [7:0] z_tempy3_G256_newbasis0;
    wire [7:0] z_cond3_G256_newbasis0;
    wire [7:0] z_negCond3_G256_newbasis0;
    wire [7:0] z_yxorb3_G256_newbasis0;
    wire [7:0] z_ny3_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond3_G256_newbasis0;
    wire [7:0] z_y3_G256_newbasis0;
    wire [7:0] z_x3_G256_newbasis0;
    wire [7:0] z_tempy4_G256_newbasis0;
    wire [7:0] z_cond4_G256_newbasis0;
    wire [7:0] z_negCond4_G256_newbasis0;
    wire [7:0] z_yxorb4_G256_newbasis0;
    wire [7:0] z_ny4_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond4_G256_newbasis0;
    wire [7:0] z_y4_G256_newbasis0;
    wire [7:0] z_x4_G256_newbasis0;
    wire [7:0] z_tempy5_G256_newbasis0;
    wire [7:0] z_cond5_G256_newbasis0;
    wire [7:0] z_negCond5_G256_newbasis0;
    wire [7:0] z_yxorb5_G256_newbasis0;
    wire [7:0] z_ny5_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond5_G256_newbasis0;
    wire [7:0] z_y5_G256_newbasis0;
    wire [7:0] z_x5_G256_newbasis0;
    wire [7:0] z_tempy6_G256_newbasis0;
    wire [7:0] z_cond6_G256_newbasis0;
    wire [7:0] z_negCond6_G256_newbasis0;
    wire [7:0] z_yxorb6_G256_newbasis0;
    wire [7:0] z_ny6_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond6_G256_newbasis0;
    wire [7:0] z_y6_G256_newbasis0;
    wire [7:0] z_x6_G256_newbasis0;
    wire [7:0] z_tempy7_G256_newbasis0;
    wire [7:0] z_cond7_G256_newbasis0;
    wire [7:0] z_negCond7_G256_newbasis0;
    wire [7:0] z_yxorb7_G256_newbasis0;
    wire [7:0] z_ny7_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond7_G256_newbasis0;
    wire [7:0] z_y7_G256_newbasis0;
    wire [7:0] z_x7_G256_newbasis0;
    wire [7:0] z_tempy8_G256_newbasis0;
    wire [7:0] z_cond8_G256_newbasis0;
    wire [7:0] z_negCond8_G256_newbasis0;
    wire [7:0] z_yxorb8_G256_newbasis0;
    wire [7:0] z_ny8_G256_newbasis0;
    wire [7:0] z_tempyIntoNegCond8_G256_newbasis0;
    wire [7:0] z_y8_G256_newbasis0;
    wire [7:0] z3285_assgn3285;
    reg [7:0] z3285_assgn32850;
    reg [7:0] z3285_assgn32851;
    reg [7:0] z3285_assgn32852;
    reg [7:0] z3285_assgn32853;
    reg [7:0] z3285_assgn32854;
    reg [7:0] z_x8_G256_newbasis0;
    wire [7:0] t3;
    wire [7:0] a0_0_G256_inv0;
    wire [7:0] a1_0_G256_inv0;
    wire [7:0] a0_G256_inv0;
    wire [7:0] a1_G256_inv0;
    wire [7:0] b0_G256_inv0;
    wire [7:0] b1_G256_inv0;
    wire [7:0] a0xorb0_G256_inv0;
    wire [7:0] a1xorb1_G256_inv0;
    wire [7:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] c0_G256_inv0;
    wire [7:0] c1_G256_inv0;
    wire [7:0] r00_G16_mul0_G256_inv0;
    wire [7:0] r10_G16_mul0_G256_inv0;
    wire [7:0] r20_G16_mul0_G256_inv0;
    wire [7:0] r30_G16_mul0_G256_inv0;
    wire [7:0] r40_G16_mul0_G256_inv0;
    wire [7:0] r50_G16_mul0_G256_inv0;
    wire [7:0] r60_G16_mul0_G256_inv0;
    wire [7:0] r70_G16_mul0_G256_inv0;
    wire [7:0] r80_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G16_mul0_G256_inv0;
    wire [7:0] a0_G16_mul0_G256_inv0;
    wire [7:0] a1_G16_mul0_G256_inv0;
    wire [7:0] b0_G16_mul0_G256_inv0;
    wire [7:0] b1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G16_mul0_G256_inv0;
    wire [7:0] c0_G16_mul0_G256_inv0;
    wire [7:0] c1_G16_mul0_G256_inv0;
    wire [7:0] d0_G16_mul0_G256_inv0;
    wire [7:0] d1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] c0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] c1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] d0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] d1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul0_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] z3583_assgn3583;
    reg [7:0] z3583_assgn35830;
    reg [7:0] z683_assgn683;
    wire [7:0] p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] z3587_assgn3587;
    reg [7:0] z3587_assgn35870;
    reg [7:0] z685_assgn685;
    wire [7:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G16_mul0_G256_inv0;
    wire [7:0] e1_G16_mul0_G256_inv0;
    wire [7:0] z3595_assgn3595;
    reg [7:0] z3595_assgn35950;
    reg [7:0] z691_assgn691;
    wire [7:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3599_assgn3599;
    reg [7:0] z3599_assgn35990;
    reg [7:0] z693_assgn693;
    wire [7:0] a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3603_assgn3603;
    reg [7:0] z3603_assgn36030;
    reg [7:0] z695_assgn695;
    wire [7:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3607_assgn3607;
    reg [7:0] z3607_assgn36070;
    reg [7:0] z697_assgn697;
    wire [7:0] a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3611_assgn3611;
    reg [7:0] z3611_assgn36110;
    reg [7:0] z699_assgn699;
    wire [7:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3615_assgn3615;
    reg [7:0] z3615_assgn36150;
    reg [7:0] z701_assgn701;
    wire [7:0] b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3627_assgn3627;
    reg [7:0] z3627_assgn36270;
    reg [7:0] z711_assgn711;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] z3631_assgn3631;
    reg [7:0] z3631_assgn36310;
    reg [7:0] z713_assgn713;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] e01_G16_mul0_G256_inv0;
    wire [7:0] e11_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] c0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] c1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] d0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] d1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul1_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] z3775_assgn3775;
    reg [7:0] z3775_assgn37750;
    reg [7:0] z855_assgn855;
    wire [7:0] p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] z3779_assgn3779;
    reg [7:0] z3779_assgn37790;
    reg [7:0] z857_assgn857;
    wire [7:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G16_mul0_G256_inv0;
    wire [7:0] p0_G16_mul0_G256_inv0;
    wire [7:0] p1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] axorb_1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] cxord_1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] c0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] c1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] u1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] b0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] d0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p0_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p1_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] b1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] d1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p2_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p3_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul2_G16_mul0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] z3927_assgn3927;
    reg [7:0] z3927_assgn39270;
    reg [7:0] z1003_assgn1003;
    wire [7:0] p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] z3931_assgn3931;
    reg [7:0] z3931_assgn39310;
    reg [7:0] z1005_assgn1005;
    wire [7:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G16_mul0_G256_inv0;
    wire [7:0] q0_G16_mul0_G256_inv0;
    wire [7:0] q1_G16_mul0_G256_inv0;
    wire [7:0] z3943_assgn3943;
    reg [7:0] z3943_assgn39430;
    reg [7:0] z1015_assgn1015;
    wire [7:0] p0ls2_G16_mul0_G256_inv0;
    wire [7:0] z3947_assgn3947;
    reg [7:0] z3947_assgn39470;
    reg [7:0] z1017_assgn1017;
    wire [7:0] p1ls2_G16_mul0_G256_inv0;
    wire [7:0] d0_G256_inv0;
    wire [7:0] d1_G256_inv0;
    wire [7:0] z3955_assgn3955;
    reg [7:0] z3955_assgn39550;
    reg [7:0] z1024_assgn1024;
    wire [7:0] c0xord0_G256_inv0;
    wire [7:0] z3959_assgn3959;
    reg [7:0] z3959_assgn39590;
    reg [7:0] z1026_assgn1026;
    wire [7:0] c1xord1_G256_inv0;
    wire [7:0] r00_G16_inv0_G256_inv0;
    wire [7:0] r10_G16_inv0_G256_inv0;
    wire [7:0] r20_G16_inv0_G256_inv0;
    wire [7:0] r30_G16_inv0_G256_inv0;
    wire [7:0] r40_G16_inv0_G256_inv0;
    wire [7:0] r50_G16_inv0_G256_inv0;
    wire [7:0] r60_G16_inv0_G256_inv0;
    wire [7:0] r70_G16_inv0_G256_inv0;
    wire [7:0] r80_G16_inv0_G256_inv0;
    wire [7:0] z3981_assgn3981;
    reg [7:0] z3981_assgn39810;
    reg [7:0] z1045_assgn1045;
    wire [7:0] a0_0_G16_inv0_G256_inv0;
    wire [7:0] z3985_assgn3985;
    reg [7:0] z3985_assgn39850;
    reg [7:0] z1047_assgn1047;
    wire [7:0] a1_0_G16_inv0_G256_inv0;
    wire [7:0] z3989_assgn3989;
    reg [7:0] z3989_assgn39890;
    reg [7:0] z1049_assgn1049;
    wire [7:0] a0_G16_inv0_G256_inv0;
    wire [7:0] z3993_assgn3993;
    reg [7:0] z3993_assgn39930;
    reg [7:0] z1051_assgn1051;
    wire [7:0] a1_G16_inv0_G256_inv0;
    wire [7:0] z3997_assgn3997;
    reg [7:0] z3997_assgn39970;
    reg [7:0] z1053_assgn1053;
    wire [7:0] b0_G16_inv0_G256_inv0;
    wire [7:0] z4001_assgn4001;
    reg [7:0] z4001_assgn40010;
    reg [7:0] z1055_assgn1055;
    wire [7:0] b1_G16_inv0_G256_inv0;
    wire [7:0] a0xorb0_G16_inv0_G256_inv0;
    wire [7:0] a1xorb1_G16_inv0_G256_inv0;
    wire [7:0] z4009_assgn4009;
    reg [7:0] z4009_assgn40090;
    reg [7:0] z1061_assgn1061;
    wire [7:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4013_assgn4013;
    reg [7:0] z4013_assgn40130;
    reg [7:0] z1063_assgn1063;
    wire [7:0] a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4017_assgn4017;
    reg [7:0] z4017_assgn40170;
    reg [7:0] z1065_assgn1065;
    wire [7:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4021_assgn4021;
    reg [7:0] z4021_assgn40210;
    reg [7:0] z1067_assgn1067;
    wire [7:0] a1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4025_assgn4025;
    reg [7:0] z4025_assgn40250;
    reg [7:0] z1069_assgn1069;
    wire [7:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4029_assgn4029;
    reg [7:0] z4029_assgn40290;
    reg [7:0] z1071_assgn1071;
    wire [7:0] b1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4033_assgn4033;
    reg [7:0] z4033_assgn40330;
    reg [7:0] z1073_assgn1073;
    wire [7:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] z4037_assgn4037;
    reg [7:0] z4037_assgn40370;
    reg [7:0] z1075_assgn1075;
    wire [7:0] b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G16_inv0_G256_inv0;
    wire [7:0] z4045_assgn4045;
    reg [7:0] z4045_assgn40450;
    reg [7:0] z1081_assgn1081;
    wire [7:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4049_assgn4049;
    reg [7:0] z4049_assgn40490;
    reg [7:0] z1083_assgn1083;
    wire [7:0] a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4053_assgn4053;
    reg [7:0] z4053_assgn40530;
    reg [7:0] z1085_assgn1085;
    wire [7:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4057_assgn4057;
    reg [7:0] z4057_assgn40570;
    reg [7:0] z1087_assgn1087;
    wire [7:0] a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4061_assgn4061;
    reg [7:0] z4061_assgn40610;
    reg [7:0] z1089_assgn1089;
    wire [7:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4065_assgn4065;
    reg [7:0] z4065_assgn40650;
    reg [7:0] z1091_assgn1091;
    wire [7:0] b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4077_assgn4077;
    reg [7:0] z4077_assgn40770;
    reg [7:0] z1101_assgn1101;
    wire [7:0] p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] z4081_assgn4081;
    reg [7:0] z4081_assgn40810;
    reg [7:0] z1103_assgn1103;
    wire [7:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] c0_G16_inv0_G256_inv0;
    wire [7:0] c1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4095_assgn4095;
    reg [7:0] z4095_assgn40950;
    reg [7:0] z1115_assgn1115;
    wire [7:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4099_assgn4099;
    reg [7:0] z4099_assgn40990;
    reg [7:0] z1117_assgn1117;
    wire [7:0] a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4103_assgn4103;
    reg [7:0] z4103_assgn41030;
    reg [7:0] z1119_assgn1119;
    wire [7:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4107_assgn4107;
    reg [7:0] z4107_assgn41070;
    reg [7:0] z1121_assgn1121;
    wire [7:0] a1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4111_assgn4111;
    reg [7:0] z4111_assgn41110;
    reg [7:0] z1123_assgn1123;
    wire [7:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4115_assgn4115;
    reg [7:0] z4115_assgn41150;
    reg [7:0] z1125_assgn1125;
    wire [7:0] b1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4119_assgn4119;
    reg [7:0] z4119_assgn41190;
    reg [7:0] z1127_assgn1127;
    wire [7:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4123_assgn4123;
    reg [7:0] z4123_assgn41230;
    reg [7:0] z1129_assgn1129;
    wire [7:0] c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4127_assgn4127;
    reg [7:0] z4127_assgn41270;
    reg [7:0] z1131_assgn1131;
    wire [7:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4131_assgn4131;
    reg [7:0] z4131_assgn41310;
    reg [7:0] z1133_assgn1133;
    wire [7:0] c1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4135_assgn4135;
    reg [7:0] z4135_assgn41350;
    reg [7:0] z1135_assgn1135;
    wire [7:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4139_assgn4139;
    reg [7:0] z4139_assgn41390;
    reg [7:0] z1137_assgn1137;
    wire [7:0] d1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4157_assgn4157;
    reg [7:0] z4157_assgn41570;
    reg [7:0] z1153_assgn1153;
    wire [7:0] u0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4161_assgn4161;
    reg [7:0] z4161_assgn41610;
    reg [7:0] z1155_assgn1155;
    wire [7:0] u1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4165_assgn4165;
    reg [7:0] z4165_assgn41650;
    reg [7:0] z1157_assgn1157;
    wire [7:0] v0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4169_assgn4169;
    reg [7:0] z4169_assgn41690;
    reg [7:0] z1159_assgn1159;
    wire [7:0] v1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4177_assgn4177;
    reg [7:0] z4177_assgn41770;
    reg [7:0] z1166_assgn1166;
    reg [7:0] p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] axorb_1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] cxord_1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4187_assgn4187;
    reg [7:0] z4187_assgn41870;
    reg [7:0] z1174_assgn1174;
    reg [7:0] p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4199_assgn4199;
    reg [7:0] z4199_assgn41990;
    reg [7:0] z1183_assgn1183;
    wire [7:0] u0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4203_assgn4203;
    reg [7:0] z4203_assgn42030;
    reg [7:0] z1185_assgn1185;
    wire [7:0] u1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4207_assgn4207;
    reg [7:0] z4207_assgn42070;
    reg [7:0] z1187_assgn1187;
    wire [7:0] v0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4211_assgn4211;
    reg [7:0] z4211_assgn42110;
    reg [7:0] z1189_assgn1189;
    wire [7:0] v1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] a0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] c0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4219_assgn4219;
    reg [7:0] z4219_assgn42190;
    reg [7:0] z1196_assgn1196;
    reg [7:0] p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] a1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] c1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc21_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4229_assgn4229;
    reg [7:0] z4229_assgn42290;
    reg [7:0] z1204_assgn1204;
    reg [7:0] p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4245_assgn4245;
    reg [7:0] z4245_assgn42450;
    reg [7:0] z1217_assgn1217;
    wire [7:0] u0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4249_assgn4249;
    reg [7:0] z4249_assgn42490;
    reg [7:0] z1219_assgn1219;
    wire [7:0] u1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4253_assgn4253;
    reg [7:0] z4253_assgn42530;
    reg [7:0] z1221_assgn1221;
    wire [7:0] v0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4257_assgn4257;
    reg [7:0] z4257_assgn42570;
    reg [7:0] z1223_assgn1223;
    wire [7:0] v1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] b0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] d0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4265_assgn4265;
    reg [7:0] z4265_assgn42650;
    reg [7:0] z1230_assgn1230;
    reg [7:0] p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] b1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [7:0] d1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p2_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p3_hpc22_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4275_assgn4275;
    reg [7:0] z4275_assgn42750;
    reg [7:0] z1238_assgn1238;
    reg [7:0] p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul3_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4285_assgn4285;
    reg [7:0] z4285_assgn42850;
    reg [7:0] z4285_assgn42851;
    reg [7:0] z4285_assgn42852;
    reg [7:0] z1245_assgn1245;
    wire [7:0] p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] z4289_assgn4289;
    reg [7:0] z4289_assgn42890;
    reg [7:0] z4289_assgn42891;
    reg [7:0] z4289_assgn42892;
    reg [7:0] z1247_assgn1247;
    wire [7:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G16_inv0_G256_inv0;
    wire [7:0] d1_G16_inv0_G256_inv0;
    wire [7:0] z4297_assgn4297;
    reg [7:0] z4297_assgn42970;
    reg [7:0] z1254_assgn1254;
    wire [7:0] c0xord0_G16_inv0_G256_inv0;
    wire [7:0] z4301_assgn4301;
    reg [7:0] z4301_assgn43010;
    reg [7:0] z1256_assgn1256;
    wire [7:0] c1xord1_G16_inv0_G256_inv0;
    wire [7:0] z4305_assgn4305;
    reg [7:0] z4305_assgn43050;
    reg [7:0] z4305_assgn43051;
    reg [7:0] z4305_assgn43052;
    reg [7:0] z1257_assgn1257;
    wire [7:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4309_assgn4309;
    reg [7:0] z4309_assgn43090;
    reg [7:0] z4309_assgn43091;
    reg [7:0] z4309_assgn43092;
    reg [7:0] z1259_assgn1259;
    wire [7:0] a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4313_assgn4313;
    reg [7:0] z4313_assgn43130;
    reg [7:0] z4313_assgn43131;
    reg [7:0] z4313_assgn43132;
    reg [7:0] z1261_assgn1261;
    wire [7:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4317_assgn4317;
    reg [7:0] z4317_assgn43170;
    reg [7:0] z4317_assgn43171;
    reg [7:0] z4317_assgn43172;
    reg [7:0] z1263_assgn1263;
    wire [7:0] a1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4321_assgn4321;
    reg [7:0] z4321_assgn43210;
    reg [7:0] z4321_assgn43211;
    reg [7:0] z4321_assgn43212;
    reg [7:0] z1265_assgn1265;
    wire [7:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4325_assgn4325;
    reg [7:0] z4325_assgn43250;
    reg [7:0] z4325_assgn43251;
    reg [7:0] z4325_assgn43252;
    reg [7:0] z1267_assgn1267;
    wire [7:0] b1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4329_assgn4329;
    reg [7:0] z4329_assgn43290;
    reg [7:0] z4329_assgn43291;
    reg [7:0] z4329_assgn43292;
    reg [7:0] z1269_assgn1269;
    wire [7:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] z4333_assgn4333;
    reg [7:0] z4333_assgn43330;
    reg [7:0] z4333_assgn43331;
    reg [7:0] z4333_assgn43332;
    reg [7:0] z1271_assgn1271;
    wire [7:0] b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] e0_G16_inv0_G256_inv0;
    wire [7:0] e1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4347_assgn4347;
    reg [7:0] z4347_assgn43470;
    reg [7:0] z4347_assgn43471;
    reg [7:0] z4347_assgn43472;
    reg [7:0] z1283_assgn1283;
    wire [7:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4351_assgn4351;
    reg [7:0] z4351_assgn43510;
    reg [7:0] z4351_assgn43511;
    reg [7:0] z4351_assgn43512;
    reg [7:0] z1285_assgn1285;
    wire [7:0] a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4355_assgn4355;
    reg [7:0] z4355_assgn43550;
    reg [7:0] z4355_assgn43551;
    reg [7:0] z4355_assgn43552;
    reg [7:0] z1287_assgn1287;
    wire [7:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4359_assgn4359;
    reg [7:0] z4359_assgn43590;
    reg [7:0] z4359_assgn43591;
    reg [7:0] z4359_assgn43592;
    reg [7:0] z1289_assgn1289;
    wire [7:0] a1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4363_assgn4363;
    reg [7:0] z4363_assgn43630;
    reg [7:0] z4363_assgn43631;
    reg [7:0] z4363_assgn43632;
    reg [7:0] z1291_assgn1291;
    wire [7:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4367_assgn4367;
    reg [7:0] z4367_assgn43670;
    reg [7:0] z4367_assgn43671;
    reg [7:0] z4367_assgn43672;
    reg [7:0] z1293_assgn1293;
    wire [7:0] b1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4371_assgn4371;
    reg [7:0] z4371_assgn43710;
    reg [7:0] z1295_assgn1295;
    wire [7:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4375_assgn4375;
    reg [7:0] z4375_assgn43750;
    reg [7:0] z1297_assgn1297;
    wire [7:0] c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4379_assgn4379;
    reg [7:0] z4379_assgn43790;
    reg [7:0] z1299_assgn1299;
    wire [7:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4383_assgn4383;
    reg [7:0] z4383_assgn43830;
    reg [7:0] z1301_assgn1301;
    wire [7:0] c1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4387_assgn4387;
    reg [7:0] z4387_assgn43870;
    reg [7:0] z1303_assgn1303;
    wire [7:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4391_assgn4391;
    reg [7:0] z4391_assgn43910;
    reg [7:0] z1305_assgn1305;
    wire [7:0] d1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4409_assgn4409;
    reg [7:0] z4409_assgn44090;
    reg [7:0] z4409_assgn44091;
    reg [7:0] z4409_assgn44092;
    reg [7:0] z1321_assgn1321;
    wire [7:0] u0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4413_assgn4413;
    reg [7:0] z4413_assgn44130;
    reg [7:0] z4413_assgn44131;
    reg [7:0] z4413_assgn44132;
    reg [7:0] z1323_assgn1323;
    wire [7:0] u1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4417_assgn4417;
    reg [7:0] z4417_assgn44170;
    reg [7:0] z1325_assgn1325;
    wire [7:0] v0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4421_assgn4421;
    reg [7:0] z4421_assgn44210;
    reg [7:0] z1327_assgn1327;
    wire [7:0] v1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4425_assgn4425;
    reg [7:0] z4425_assgn44250;
    reg [7:0] z1329_assgn1329;
    wire [7:0] p0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4429_assgn4429;
    reg [7:0] z4429_assgn44290;
    reg [7:0] z1331_assgn1331;
    wire [7:0] p1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4437_assgn4437;
    reg [7:0] z4437_assgn44370;
    reg [7:0] z1337_assgn1337;
    wire [7:0] p2_hpc20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4441_assgn4441;
    reg [7:0] z4441_assgn44410;
    reg [7:0] z1339_assgn1339;
    wire [7:0] p3_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4455_assgn4455;
    reg [7:0] z4455_assgn44550;
    reg [7:0] z4455_assgn44551;
    reg [7:0] z4455_assgn44552;
    reg [7:0] z1351_assgn1351;
    wire [7:0] u0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4459_assgn4459;
    reg [7:0] z4459_assgn44590;
    reg [7:0] z4459_assgn44591;
    reg [7:0] z4459_assgn44592;
    reg [7:0] z1353_assgn1353;
    wire [7:0] u1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4463_assgn4463;
    reg [7:0] z4463_assgn44630;
    reg [7:0] z1355_assgn1355;
    wire [7:0] v0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4467_assgn4467;
    reg [7:0] z4467_assgn44670;
    reg [7:0] z1357_assgn1357;
    wire [7:0] v1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4471_assgn4471;
    reg [7:0] z4471_assgn44710;
    reg [7:0] z1359_assgn1359;
    wire [7:0] p0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4475_assgn4475;
    reg [7:0] z4475_assgn44750;
    reg [7:0] z1361_assgn1361;
    wire [7:0] p1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4483_assgn4483;
    reg [7:0] z4483_assgn44830;
    reg [7:0] z1367_assgn1367;
    wire [7:0] p2_hpc21_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4487_assgn4487;
    reg [7:0] z4487_assgn44870;
    reg [7:0] z1369_assgn1369;
    wire [7:0] p3_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4505_assgn4505;
    reg [7:0] z4505_assgn45050;
    reg [7:0] z4505_assgn45051;
    reg [7:0] z4505_assgn45052;
    reg [7:0] z1385_assgn1385;
    wire [7:0] u0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4509_assgn4509;
    reg [7:0] z4509_assgn45090;
    reg [7:0] z4509_assgn45091;
    reg [7:0] z4509_assgn45092;
    reg [7:0] z1387_assgn1387;
    wire [7:0] u1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4513_assgn4513;
    reg [7:0] z4513_assgn45130;
    reg [7:0] z1389_assgn1389;
    wire [7:0] v0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4517_assgn4517;
    reg [7:0] z4517_assgn45170;
    reg [7:0] z1391_assgn1391;
    wire [7:0] v1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4521_assgn4521;
    reg [7:0] z4521_assgn45210;
    reg [7:0] z1393_assgn1393;
    wire [7:0] p0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4525_assgn4525;
    reg [7:0] z4525_assgn45250;
    reg [7:0] z1395_assgn1395;
    wire [7:0] p1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4533_assgn4533;
    reg [7:0] z4533_assgn45330;
    reg [7:0] z1401_assgn1401;
    wire [7:0] p2_hpc22_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4537_assgn4537;
    reg [7:0] z4537_assgn45370;
    reg [7:0] z1403_assgn1403;
    wire [7:0] p3_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul4_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4549_assgn4549;
    reg [7:0] z4549_assgn45490;
    reg [7:0] z4549_assgn45491;
    reg [7:0] z4549_assgn45492;
    reg [7:0] z4549_assgn45493;
    reg [7:0] z1413_assgn1413;
    wire [7:0] p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] z4553_assgn4553;
    reg [7:0] z4553_assgn45530;
    reg [7:0] z4553_assgn45531;
    reg [7:0] z4553_assgn45532;
    reg [7:0] z4553_assgn45533;
    reg [7:0] z1415_assgn1415;
    wire [7:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G16_inv0_G256_inv0;
    wire [7:0] p1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4567_assgn4567;
    reg [7:0] z4567_assgn45670;
    reg [7:0] z4567_assgn45671;
    reg [7:0] z4567_assgn45672;
    reg [7:0] z1427_assgn1427;
    wire [7:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4571_assgn4571;
    reg [7:0] z4571_assgn45710;
    reg [7:0] z4571_assgn45711;
    reg [7:0] z4571_assgn45712;
    reg [7:0] z1429_assgn1429;
    wire [7:0] a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4575_assgn4575;
    reg [7:0] z4575_assgn45750;
    reg [7:0] z4575_assgn45751;
    reg [7:0] z4575_assgn45752;
    reg [7:0] z1431_assgn1431;
    wire [7:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4579_assgn4579;
    reg [7:0] z4579_assgn45790;
    reg [7:0] z4579_assgn45791;
    reg [7:0] z4579_assgn45792;
    reg [7:0] z1433_assgn1433;
    wire [7:0] a1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4583_assgn4583;
    reg [7:0] z4583_assgn45830;
    reg [7:0] z4583_assgn45831;
    reg [7:0] z4583_assgn45832;
    reg [7:0] z1435_assgn1435;
    wire [7:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4587_assgn4587;
    reg [7:0] z4587_assgn45870;
    reg [7:0] z4587_assgn45871;
    reg [7:0] z4587_assgn45872;
    reg [7:0] z1437_assgn1437;
    wire [7:0] b1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4591_assgn4591;
    reg [7:0] z4591_assgn45910;
    reg [7:0] z1439_assgn1439;
    wire [7:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4595_assgn4595;
    reg [7:0] z4595_assgn45950;
    reg [7:0] z1441_assgn1441;
    wire [7:0] c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4599_assgn4599;
    reg [7:0] z4599_assgn45990;
    reg [7:0] z1443_assgn1443;
    wire [7:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4603_assgn4603;
    reg [7:0] z4603_assgn46030;
    reg [7:0] z1445_assgn1445;
    wire [7:0] c1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4607_assgn4607;
    reg [7:0] z4607_assgn46070;
    reg [7:0] z1447_assgn1447;
    wire [7:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4611_assgn4611;
    reg [7:0] z4611_assgn46110;
    reg [7:0] z1449_assgn1449;
    wire [7:0] d1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4629_assgn4629;
    reg [7:0] z4629_assgn46290;
    reg [7:0] z4629_assgn46291;
    reg [7:0] z4629_assgn46292;
    reg [7:0] z1465_assgn1465;
    wire [7:0] u0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4633_assgn4633;
    reg [7:0] z4633_assgn46330;
    reg [7:0] z4633_assgn46331;
    reg [7:0] z4633_assgn46332;
    reg [7:0] z1467_assgn1467;
    wire [7:0] u1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4637_assgn4637;
    reg [7:0] z4637_assgn46370;
    reg [7:0] z1469_assgn1469;
    wire [7:0] v0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4641_assgn4641;
    reg [7:0] z4641_assgn46410;
    reg [7:0] z1471_assgn1471;
    wire [7:0] v1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4645_assgn4645;
    reg [7:0] z4645_assgn46450;
    reg [7:0] z1473_assgn1473;
    wire [7:0] p0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4649_assgn4649;
    reg [7:0] z4649_assgn46490;
    reg [7:0] z1475_assgn1475;
    wire [7:0] p1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] e0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4657_assgn4657;
    reg [7:0] z4657_assgn46570;
    reg [7:0] z1481_assgn1481;
    wire [7:0] p2_hpc20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4661_assgn4661;
    reg [7:0] z4661_assgn46610;
    reg [7:0] z1483_assgn1483;
    wire [7:0] p3_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] e1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4675_assgn4675;
    reg [7:0] z4675_assgn46750;
    reg [7:0] z4675_assgn46751;
    reg [7:0] z4675_assgn46752;
    reg [7:0] z1495_assgn1495;
    wire [7:0] u0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4679_assgn4679;
    reg [7:0] z4679_assgn46790;
    reg [7:0] z4679_assgn46791;
    reg [7:0] z4679_assgn46792;
    reg [7:0] z1497_assgn1497;
    wire [7:0] u1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4683_assgn4683;
    reg [7:0] z4683_assgn46830;
    reg [7:0] z1499_assgn1499;
    wire [7:0] v0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4687_assgn4687;
    reg [7:0] z4687_assgn46870;
    reg [7:0] z1501_assgn1501;
    wire [7:0] v1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4691_assgn4691;
    reg [7:0] z4691_assgn46910;
    reg [7:0] z1503_assgn1503;
    wire [7:0] p0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4695_assgn4695;
    reg [7:0] z4695_assgn46950;
    reg [7:0] z1505_assgn1505;
    wire [7:0] p1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4703_assgn4703;
    reg [7:0] z4703_assgn47030;
    reg [7:0] z1511_assgn1511;
    wire [7:0] p2_hpc21_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4707_assgn4707;
    reg [7:0] z4707_assgn47070;
    reg [7:0] z1513_assgn1513;
    wire [7:0] p3_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4725_assgn4725;
    reg [7:0] z4725_assgn47250;
    reg [7:0] z4725_assgn47251;
    reg [7:0] z4725_assgn47252;
    reg [7:0] z1529_assgn1529;
    wire [7:0] u0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4729_assgn4729;
    reg [7:0] z4729_assgn47290;
    reg [7:0] z4729_assgn47291;
    reg [7:0] z4729_assgn47292;
    reg [7:0] z1531_assgn1531;
    wire [7:0] u1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4733_assgn4733;
    reg [7:0] z4733_assgn47330;
    reg [7:0] z1533_assgn1533;
    wire [7:0] v0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4737_assgn4737;
    reg [7:0] z4737_assgn47370;
    reg [7:0] z1535_assgn1535;
    wire [7:0] v1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4741_assgn4741;
    reg [7:0] z4741_assgn47410;
    reg [7:0] z1537_assgn1537;
    wire [7:0] p0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4745_assgn4745;
    reg [7:0] z4745_assgn47450;
    reg [7:0] z1539_assgn1539;
    wire [7:0] p1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4753_assgn4753;
    reg [7:0] z4753_assgn47530;
    reg [7:0] z1545_assgn1545;
    wire [7:0] p2_hpc22_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4757_assgn4757;
    reg [7:0] z4757_assgn47570;
    reg [7:0] z1547_assgn1547;
    wire [7:0] p3_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul5_G16_inv0_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4769_assgn4769;
    reg [7:0] z4769_assgn47690;
    reg [7:0] z4769_assgn47691;
    reg [7:0] z4769_assgn47692;
    reg [7:0] z4769_assgn47693;
    reg [7:0] z1557_assgn1557;
    wire [7:0] p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] z4773_assgn4773;
    reg [7:0] z4773_assgn47730;
    reg [7:0] z4773_assgn47731;
    reg [7:0] z4773_assgn47732;
    reg [7:0] z4773_assgn47733;
    reg [7:0] z1559_assgn1559;
    wire [7:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G16_inv0_G256_inv0;
    wire [7:0] q1_G16_inv0_G256_inv0;
    wire [7:0] z4781_assgn4781;
    reg [7:0] z4781_assgn47810;
    reg [7:0] z4781_assgn47811;
    reg [7:0] z4781_assgn47812;
    reg [7:0] z4781_assgn47813;
    reg [7:0] z1565_assgn1565;
    wire [7:0] p0ls2_G16_inv0_G256_inv0;
    wire [7:0] z4785_assgn4785;
    reg [7:0] z4785_assgn47850;
    reg [7:0] z4785_assgn47851;
    reg [7:0] z4785_assgn47852;
    reg [7:0] z4785_assgn47853;
    reg [7:0] z1567_assgn1567;
    wire [7:0] p1ls2_G16_inv0_G256_inv0;
    wire [7:0] e0_G256_inv0;
    wire [7:0] e1_G256_inv0;
    wire [7:0] r00_G16_mul1_G256_inv0;
    wire [7:0] r10_G16_mul1_G256_inv0;
    wire [7:0] r20_G16_mul1_G256_inv0;
    wire [7:0] r30_G16_mul1_G256_inv0;
    wire [7:0] r40_G16_mul1_G256_inv0;
    wire [7:0] r50_G16_mul1_G256_inv0;
    wire [7:0] r60_G16_mul1_G256_inv0;
    wire [7:0] r70_G16_mul1_G256_inv0;
    wire [7:0] r80_G16_mul1_G256_inv0;
    wire [7:0] z4811_assgn4811;
    reg [7:0] z4811_assgn48110;
    reg [7:0] z4811_assgn48111;
    reg [7:0] z4811_assgn48112;
    reg [7:0] z4811_assgn48113;
    reg [7:0] z1591_assgn1591;
    wire [7:0] a0_0_G16_mul1_G256_inv0;
    wire [7:0] z4815_assgn4815;
    reg [7:0] z4815_assgn48150;
    reg [7:0] z4815_assgn48151;
    reg [7:0] z4815_assgn48152;
    reg [7:0] z4815_assgn48153;
    reg [7:0] z1593_assgn1593;
    wire [7:0] a1_0_G16_mul1_G256_inv0;
    wire [7:0] z4819_assgn4819;
    reg [7:0] z4819_assgn48190;
    reg [7:0] z4819_assgn48191;
    reg [7:0] z4819_assgn48192;
    reg [7:0] z4819_assgn48193;
    reg [7:0] z1595_assgn1595;
    wire [7:0] a0_G16_mul1_G256_inv0;
    wire [7:0] z4823_assgn4823;
    reg [7:0] z4823_assgn48230;
    reg [7:0] z4823_assgn48231;
    reg [7:0] z4823_assgn48232;
    reg [7:0] z4823_assgn48233;
    reg [7:0] z1597_assgn1597;
    wire [7:0] a1_G16_mul1_G256_inv0;
    wire [7:0] z4827_assgn4827;
    reg [7:0] z4827_assgn48270;
    reg [7:0] z4827_assgn48271;
    reg [7:0] z4827_assgn48272;
    reg [7:0] z4827_assgn48273;
    reg [7:0] z1599_assgn1599;
    wire [7:0] b0_G16_mul1_G256_inv0;
    wire [7:0] z4831_assgn4831;
    reg [7:0] z4831_assgn48310;
    reg [7:0] z4831_assgn48311;
    reg [7:0] z4831_assgn48312;
    reg [7:0] z4831_assgn48313;
    reg [7:0] z1601_assgn1601;
    wire [7:0] b1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G16_mul1_G256_inv0;
    wire [7:0] c0_G16_mul1_G256_inv0;
    wire [7:0] c1_G16_mul1_G256_inv0;
    wire [7:0] d0_G16_mul1_G256_inv0;
    wire [7:0] d1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4861_assgn4861;
    reg [7:0] z4861_assgn48610;
    reg [7:0] z4861_assgn48611;
    reg [7:0] z4861_assgn48612;
    reg [7:0] z4861_assgn48613;
    reg [7:0] z1629_assgn1629;
    wire [7:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4865_assgn4865;
    reg [7:0] z4865_assgn48650;
    reg [7:0] z4865_assgn48651;
    reg [7:0] z4865_assgn48652;
    reg [7:0] z4865_assgn48653;
    reg [7:0] z1631_assgn1631;
    wire [7:0] a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4869_assgn4869;
    reg [7:0] z4869_assgn48690;
    reg [7:0] z4869_assgn48691;
    reg [7:0] z4869_assgn48692;
    reg [7:0] z4869_assgn48693;
    reg [7:0] z1633_assgn1633;
    wire [7:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4873_assgn4873;
    reg [7:0] z4873_assgn48730;
    reg [7:0] z4873_assgn48731;
    reg [7:0] z4873_assgn48732;
    reg [7:0] z4873_assgn48733;
    reg [7:0] z1635_assgn1635;
    wire [7:0] a1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4877_assgn4877;
    reg [7:0] z4877_assgn48770;
    reg [7:0] z4877_assgn48771;
    reg [7:0] z4877_assgn48772;
    reg [7:0] z4877_assgn48773;
    reg [7:0] z1637_assgn1637;
    wire [7:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4881_assgn4881;
    reg [7:0] z4881_assgn48810;
    reg [7:0] z4881_assgn48811;
    reg [7:0] z4881_assgn48812;
    reg [7:0] z4881_assgn48813;
    reg [7:0] z1639_assgn1639;
    wire [7:0] b1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4911_assgn4911;
    reg [7:0] z4911_assgn49110;
    reg [7:0] z4911_assgn49111;
    reg [7:0] z4911_assgn49112;
    reg [7:0] z4911_assgn49113;
    reg [7:0] z1667_assgn1667;
    wire [7:0] u0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4915_assgn4915;
    reg [7:0] z4915_assgn49150;
    reg [7:0] z4915_assgn49151;
    reg [7:0] z4915_assgn49152;
    reg [7:0] z4915_assgn49153;
    reg [7:0] z1669_assgn1669;
    wire [7:0] u1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4923_assgn4923;
    reg [7:0] z4923_assgn49230;
    reg [7:0] z4923_assgn49231;
    reg [7:0] z4923_assgn49232;
    reg [7:0] z4923_assgn49233;
    reg [7:0] z1675_assgn1675;
    wire [7:0] p0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4927_assgn4927;
    reg [7:0] z4927_assgn49270;
    reg [7:0] z4927_assgn49271;
    reg [7:0] z4927_assgn49272;
    reg [7:0] z4927_assgn49273;
    reg [7:0] z1677_assgn1677;
    wire [7:0] p1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4935_assgn4935;
    reg [7:0] z4935_assgn49350;
    reg [7:0] z4935_assgn49351;
    reg [7:0] z4935_assgn49352;
    reg [7:0] z4935_assgn49353;
    reg [7:0] z1683_assgn1683;
    wire [7:0] p2_hpc20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4939_assgn4939;
    reg [7:0] z4939_assgn49390;
    reg [7:0] z4939_assgn49391;
    reg [7:0] z4939_assgn49392;
    reg [7:0] z4939_assgn49393;
    reg [7:0] z1685_assgn1685;
    wire [7:0] p3_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4953_assgn4953;
    reg [7:0] z4953_assgn49530;
    reg [7:0] z4953_assgn49531;
    reg [7:0] z4953_assgn49532;
    reg [7:0] z4953_assgn49533;
    reg [7:0] z1697_assgn1697;
    wire [7:0] u0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4957_assgn4957;
    reg [7:0] z4957_assgn49570;
    reg [7:0] z4957_assgn49571;
    reg [7:0] z4957_assgn49572;
    reg [7:0] z4957_assgn49573;
    reg [7:0] z1699_assgn1699;
    wire [7:0] u1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4965_assgn4965;
    reg [7:0] z4965_assgn49650;
    reg [7:0] z4965_assgn49651;
    reg [7:0] z4965_assgn49652;
    reg [7:0] z4965_assgn49653;
    reg [7:0] z1705_assgn1705;
    wire [7:0] p0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4969_assgn4969;
    reg [7:0] z4969_assgn49690;
    reg [7:0] z4969_assgn49691;
    reg [7:0] z4969_assgn49692;
    reg [7:0] z4969_assgn49693;
    reg [7:0] z1707_assgn1707;
    wire [7:0] p1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4977_assgn4977;
    reg [7:0] z4977_assgn49770;
    reg [7:0] z4977_assgn49771;
    reg [7:0] z4977_assgn49772;
    reg [7:0] z4977_assgn49773;
    reg [7:0] z1713_assgn1713;
    wire [7:0] p2_hpc21_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4981_assgn4981;
    reg [7:0] z4981_assgn49810;
    reg [7:0] z4981_assgn49811;
    reg [7:0] z4981_assgn49812;
    reg [7:0] z4981_assgn49813;
    reg [7:0] z1715_assgn1715;
    wire [7:0] p3_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z4999_assgn4999;
    reg [7:0] z4999_assgn49990;
    reg [7:0] z4999_assgn49991;
    reg [7:0] z4999_assgn49992;
    reg [7:0] z4999_assgn49993;
    reg [7:0] z1731_assgn1731;
    wire [7:0] u0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5003_assgn5003;
    reg [7:0] z5003_assgn50030;
    reg [7:0] z5003_assgn50031;
    reg [7:0] z5003_assgn50032;
    reg [7:0] z5003_assgn50033;
    reg [7:0] z1733_assgn1733;
    wire [7:0] u1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5011_assgn5011;
    reg [7:0] z5011_assgn50110;
    reg [7:0] z5011_assgn50111;
    reg [7:0] z5011_assgn50112;
    reg [7:0] z5011_assgn50113;
    reg [7:0] z1739_assgn1739;
    wire [7:0] p0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5015_assgn5015;
    reg [7:0] z5015_assgn50150;
    reg [7:0] z5015_assgn50151;
    reg [7:0] z5015_assgn50152;
    reg [7:0] z5015_assgn50153;
    reg [7:0] z1741_assgn1741;
    wire [7:0] p1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5023_assgn5023;
    reg [7:0] z5023_assgn50230;
    reg [7:0] z5023_assgn50231;
    reg [7:0] z5023_assgn50232;
    reg [7:0] z5023_assgn50233;
    reg [7:0] z1747_assgn1747;
    wire [7:0] p2_hpc22_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5027_assgn5027;
    reg [7:0] z5027_assgn50270;
    reg [7:0] z5027_assgn50271;
    reg [7:0] z5027_assgn50272;
    reg [7:0] z5027_assgn50273;
    reg [7:0] z1749_assgn1749;
    wire [7:0] p3_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul0_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5039_assgn5039;
    reg [7:0] z5039_assgn50390;
    reg [7:0] z5039_assgn50391;
    reg [7:0] z5039_assgn50392;
    reg [7:0] z5039_assgn50393;
    reg [7:0] z5039_assgn50394;
    reg [7:0] z1759_assgn1759;
    wire [7:0] p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] z5043_assgn5043;
    reg [7:0] z5043_assgn50430;
    reg [7:0] z5043_assgn50431;
    reg [7:0] z5043_assgn50432;
    reg [7:0] z5043_assgn50433;
    reg [7:0] z5043_assgn50434;
    reg [7:0] z1761_assgn1761;
    wire [7:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G16_mul1_G256_inv0;
    wire [7:0] e1_G16_mul1_G256_inv0;
    wire [7:0] z5051_assgn5051;
    reg [7:0] z5051_assgn50510;
    reg [7:0] z5051_assgn50511;
    reg [7:0] z5051_assgn50512;
    reg [7:0] z5051_assgn50513;
    reg [7:0] z5051_assgn50514;
    reg [7:0] z1767_assgn1767;
    wire [7:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5055_assgn5055;
    reg [7:0] z5055_assgn50550;
    reg [7:0] z5055_assgn50551;
    reg [7:0] z5055_assgn50552;
    reg [7:0] z5055_assgn50553;
    reg [7:0] z5055_assgn50554;
    reg [7:0] z1769_assgn1769;
    wire [7:0] a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5059_assgn5059;
    reg [7:0] z5059_assgn50590;
    reg [7:0] z5059_assgn50591;
    reg [7:0] z5059_assgn50592;
    reg [7:0] z5059_assgn50593;
    reg [7:0] z5059_assgn50594;
    reg [7:0] z1771_assgn1771;
    wire [7:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5063_assgn5063;
    reg [7:0] z5063_assgn50630;
    reg [7:0] z5063_assgn50631;
    reg [7:0] z5063_assgn50632;
    reg [7:0] z5063_assgn50633;
    reg [7:0] z5063_assgn50634;
    reg [7:0] z1773_assgn1773;
    wire [7:0] a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5067_assgn5067;
    reg [7:0] z5067_assgn50670;
    reg [7:0] z5067_assgn50671;
    reg [7:0] z5067_assgn50672;
    reg [7:0] z5067_assgn50673;
    reg [7:0] z5067_assgn50674;
    reg [7:0] z1775_assgn1775;
    wire [7:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5071_assgn5071;
    reg [7:0] z5071_assgn50710;
    reg [7:0] z5071_assgn50711;
    reg [7:0] z5071_assgn50712;
    reg [7:0] z5071_assgn50713;
    reg [7:0] z5071_assgn50714;
    reg [7:0] z1777_assgn1777;
    wire [7:0] b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5083_assgn5083;
    reg [7:0] z5083_assgn50830;
    reg [7:0] z5083_assgn50831;
    reg [7:0] z5083_assgn50832;
    reg [7:0] z5083_assgn50833;
    reg [7:0] z5083_assgn50834;
    reg [7:0] z1787_assgn1787;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] z5087_assgn5087;
    reg [7:0] z5087_assgn50870;
    reg [7:0] z5087_assgn50871;
    reg [7:0] z5087_assgn50872;
    reg [7:0] z5087_assgn50873;
    reg [7:0] z5087_assgn50874;
    reg [7:0] z1789_assgn1789;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] e01_G16_mul1_G256_inv0;
    wire [7:0] e11_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5101_assgn5101;
    reg [7:0] z5101_assgn51010;
    reg [7:0] z5101_assgn51011;
    reg [7:0] z5101_assgn51012;
    reg [7:0] z5101_assgn51013;
    reg [7:0] z1801_assgn1801;
    wire [7:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5105_assgn5105;
    reg [7:0] z5105_assgn51050;
    reg [7:0] z5105_assgn51051;
    reg [7:0] z5105_assgn51052;
    reg [7:0] z5105_assgn51053;
    reg [7:0] z1803_assgn1803;
    wire [7:0] a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5109_assgn5109;
    reg [7:0] z5109_assgn51090;
    reg [7:0] z5109_assgn51091;
    reg [7:0] z5109_assgn51092;
    reg [7:0] z5109_assgn51093;
    reg [7:0] z1805_assgn1805;
    wire [7:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5113_assgn5113;
    reg [7:0] z5113_assgn51130;
    reg [7:0] z5113_assgn51131;
    reg [7:0] z5113_assgn51132;
    reg [7:0] z5113_assgn51133;
    reg [7:0] z1807_assgn1807;
    wire [7:0] a1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5117_assgn5117;
    reg [7:0] z5117_assgn51170;
    reg [7:0] z5117_assgn51171;
    reg [7:0] z5117_assgn51172;
    reg [7:0] z5117_assgn51173;
    reg [7:0] z1809_assgn1809;
    wire [7:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5121_assgn5121;
    reg [7:0] z5121_assgn51210;
    reg [7:0] z5121_assgn51211;
    reg [7:0] z5121_assgn51212;
    reg [7:0] z5121_assgn51213;
    reg [7:0] z1811_assgn1811;
    wire [7:0] b1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5151_assgn5151;
    reg [7:0] z5151_assgn51510;
    reg [7:0] z5151_assgn51511;
    reg [7:0] z5151_assgn51512;
    reg [7:0] z5151_assgn51513;
    reg [7:0] z1839_assgn1839;
    wire [7:0] u0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5155_assgn5155;
    reg [7:0] z5155_assgn51550;
    reg [7:0] z5155_assgn51551;
    reg [7:0] z5155_assgn51552;
    reg [7:0] z5155_assgn51553;
    reg [7:0] z1841_assgn1841;
    wire [7:0] u1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5163_assgn5163;
    reg [7:0] z5163_assgn51630;
    reg [7:0] z5163_assgn51631;
    reg [7:0] z5163_assgn51632;
    reg [7:0] z5163_assgn51633;
    reg [7:0] z1847_assgn1847;
    wire [7:0] p0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5167_assgn5167;
    reg [7:0] z5167_assgn51670;
    reg [7:0] z5167_assgn51671;
    reg [7:0] z5167_assgn51672;
    reg [7:0] z5167_assgn51673;
    reg [7:0] z1849_assgn1849;
    wire [7:0] p1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5175_assgn5175;
    reg [7:0] z5175_assgn51750;
    reg [7:0] z5175_assgn51751;
    reg [7:0] z5175_assgn51752;
    reg [7:0] z5175_assgn51753;
    reg [7:0] z1855_assgn1855;
    wire [7:0] p2_hpc20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5179_assgn5179;
    reg [7:0] z5179_assgn51790;
    reg [7:0] z5179_assgn51791;
    reg [7:0] z5179_assgn51792;
    reg [7:0] z5179_assgn51793;
    reg [7:0] z1857_assgn1857;
    wire [7:0] p3_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5193_assgn5193;
    reg [7:0] z5193_assgn51930;
    reg [7:0] z5193_assgn51931;
    reg [7:0] z5193_assgn51932;
    reg [7:0] z5193_assgn51933;
    reg [7:0] z1869_assgn1869;
    wire [7:0] u0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5197_assgn5197;
    reg [7:0] z5197_assgn51970;
    reg [7:0] z5197_assgn51971;
    reg [7:0] z5197_assgn51972;
    reg [7:0] z5197_assgn51973;
    reg [7:0] z1871_assgn1871;
    wire [7:0] u1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5205_assgn5205;
    reg [7:0] z5205_assgn52050;
    reg [7:0] z5205_assgn52051;
    reg [7:0] z5205_assgn52052;
    reg [7:0] z5205_assgn52053;
    reg [7:0] z1877_assgn1877;
    wire [7:0] p0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5209_assgn5209;
    reg [7:0] z5209_assgn52090;
    reg [7:0] z5209_assgn52091;
    reg [7:0] z5209_assgn52092;
    reg [7:0] z5209_assgn52093;
    reg [7:0] z1879_assgn1879;
    wire [7:0] p1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5217_assgn5217;
    reg [7:0] z5217_assgn52170;
    reg [7:0] z5217_assgn52171;
    reg [7:0] z5217_assgn52172;
    reg [7:0] z5217_assgn52173;
    reg [7:0] z1885_assgn1885;
    wire [7:0] p2_hpc21_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5221_assgn5221;
    reg [7:0] z5221_assgn52210;
    reg [7:0] z5221_assgn52211;
    reg [7:0] z5221_assgn52212;
    reg [7:0] z5221_assgn52213;
    reg [7:0] z1887_assgn1887;
    wire [7:0] p3_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5239_assgn5239;
    reg [7:0] z5239_assgn52390;
    reg [7:0] z5239_assgn52391;
    reg [7:0] z5239_assgn52392;
    reg [7:0] z5239_assgn52393;
    reg [7:0] z1903_assgn1903;
    wire [7:0] u0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5243_assgn5243;
    reg [7:0] z5243_assgn52430;
    reg [7:0] z5243_assgn52431;
    reg [7:0] z5243_assgn52432;
    reg [7:0] z5243_assgn52433;
    reg [7:0] z1905_assgn1905;
    wire [7:0] u1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5251_assgn5251;
    reg [7:0] z5251_assgn52510;
    reg [7:0] z5251_assgn52511;
    reg [7:0] z5251_assgn52512;
    reg [7:0] z5251_assgn52513;
    reg [7:0] z1911_assgn1911;
    wire [7:0] p0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5255_assgn5255;
    reg [7:0] z5255_assgn52550;
    reg [7:0] z5255_assgn52551;
    reg [7:0] z5255_assgn52552;
    reg [7:0] z5255_assgn52553;
    reg [7:0] z1913_assgn1913;
    wire [7:0] p1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5263_assgn5263;
    reg [7:0] z5263_assgn52630;
    reg [7:0] z5263_assgn52631;
    reg [7:0] z5263_assgn52632;
    reg [7:0] z5263_assgn52633;
    reg [7:0] z1919_assgn1919;
    wire [7:0] p2_hpc22_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5267_assgn5267;
    reg [7:0] z5267_assgn52670;
    reg [7:0] z5267_assgn52671;
    reg [7:0] z5267_assgn52672;
    reg [7:0] z5267_assgn52673;
    reg [7:0] z1921_assgn1921;
    wire [7:0] p3_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul1_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5279_assgn5279;
    reg [7:0] z5279_assgn52790;
    reg [7:0] z5279_assgn52791;
    reg [7:0] z5279_assgn52792;
    reg [7:0] z5279_assgn52793;
    reg [7:0] z5279_assgn52794;
    reg [7:0] z1931_assgn1931;
    wire [7:0] p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] z5283_assgn5283;
    reg [7:0] z5283_assgn52830;
    reg [7:0] z5283_assgn52831;
    reg [7:0] z5283_assgn52832;
    reg [7:0] z5283_assgn52833;
    reg [7:0] z5283_assgn52834;
    reg [7:0] z1933_assgn1933;
    wire [7:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G16_mul1_G256_inv0;
    wire [7:0] p0_G16_mul1_G256_inv0;
    wire [7:0] p1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5301_assgn5301;
    reg [7:0] z5301_assgn53010;
    reg [7:0] z5301_assgn53011;
    reg [7:0] z5301_assgn53012;
    reg [7:0] z5301_assgn53013;
    reg [7:0] z1949_assgn1949;
    wire [7:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5305_assgn5305;
    reg [7:0] z5305_assgn53050;
    reg [7:0] z5305_assgn53051;
    reg [7:0] z5305_assgn53052;
    reg [7:0] z5305_assgn53053;
    reg [7:0] z1951_assgn1951;
    wire [7:0] a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5309_assgn5309;
    reg [7:0] z5309_assgn53090;
    reg [7:0] z5309_assgn53091;
    reg [7:0] z5309_assgn53092;
    reg [7:0] z5309_assgn53093;
    reg [7:0] z1953_assgn1953;
    wire [7:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5313_assgn5313;
    reg [7:0] z5313_assgn53130;
    reg [7:0] z5313_assgn53131;
    reg [7:0] z5313_assgn53132;
    reg [7:0] z5313_assgn53133;
    reg [7:0] z1955_assgn1955;
    wire [7:0] a1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5317_assgn5317;
    reg [7:0] z5317_assgn53170;
    reg [7:0] z5317_assgn53171;
    reg [7:0] z5317_assgn53172;
    reg [7:0] z5317_assgn53173;
    reg [7:0] z1957_assgn1957;
    wire [7:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5321_assgn5321;
    reg [7:0] z5321_assgn53210;
    reg [7:0] z5321_assgn53211;
    reg [7:0] z5321_assgn53212;
    reg [7:0] z5321_assgn53213;
    reg [7:0] z1959_assgn1959;
    wire [7:0] b1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5351_assgn5351;
    reg [7:0] z5351_assgn53510;
    reg [7:0] z5351_assgn53511;
    reg [7:0] z5351_assgn53512;
    reg [7:0] z5351_assgn53513;
    reg [7:0] z1987_assgn1987;
    wire [7:0] u0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5355_assgn5355;
    reg [7:0] z5355_assgn53550;
    reg [7:0] z5355_assgn53551;
    reg [7:0] z5355_assgn53552;
    reg [7:0] z5355_assgn53553;
    reg [7:0] z1989_assgn1989;
    wire [7:0] u1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5363_assgn5363;
    reg [7:0] z5363_assgn53630;
    reg [7:0] z5363_assgn53631;
    reg [7:0] z5363_assgn53632;
    reg [7:0] z5363_assgn53633;
    reg [7:0] z1995_assgn1995;
    wire [7:0] p0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5367_assgn5367;
    reg [7:0] z5367_assgn53670;
    reg [7:0] z5367_assgn53671;
    reg [7:0] z5367_assgn53672;
    reg [7:0] z5367_assgn53673;
    reg [7:0] z1997_assgn1997;
    wire [7:0] p1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5375_assgn5375;
    reg [7:0] z5375_assgn53750;
    reg [7:0] z5375_assgn53751;
    reg [7:0] z5375_assgn53752;
    reg [7:0] z5375_assgn53753;
    reg [7:0] z2003_assgn2003;
    wire [7:0] p2_hpc20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5379_assgn5379;
    reg [7:0] z5379_assgn53790;
    reg [7:0] z5379_assgn53791;
    reg [7:0] z5379_assgn53792;
    reg [7:0] z5379_assgn53793;
    reg [7:0] z2005_assgn2005;
    wire [7:0] p3_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5393_assgn5393;
    reg [7:0] z5393_assgn53930;
    reg [7:0] z5393_assgn53931;
    reg [7:0] z5393_assgn53932;
    reg [7:0] z5393_assgn53933;
    reg [7:0] z2017_assgn2017;
    wire [7:0] u0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5397_assgn5397;
    reg [7:0] z5397_assgn53970;
    reg [7:0] z5397_assgn53971;
    reg [7:0] z5397_assgn53972;
    reg [7:0] z5397_assgn53973;
    reg [7:0] z2019_assgn2019;
    wire [7:0] u1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5405_assgn5405;
    reg [7:0] z5405_assgn54050;
    reg [7:0] z5405_assgn54051;
    reg [7:0] z5405_assgn54052;
    reg [7:0] z5405_assgn54053;
    reg [7:0] z2025_assgn2025;
    wire [7:0] p0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5409_assgn5409;
    reg [7:0] z5409_assgn54090;
    reg [7:0] z5409_assgn54091;
    reg [7:0] z5409_assgn54092;
    reg [7:0] z5409_assgn54093;
    reg [7:0] z2027_assgn2027;
    wire [7:0] p1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5417_assgn5417;
    reg [7:0] z5417_assgn54170;
    reg [7:0] z5417_assgn54171;
    reg [7:0] z5417_assgn54172;
    reg [7:0] z5417_assgn54173;
    reg [7:0] z2033_assgn2033;
    wire [7:0] p2_hpc21_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5421_assgn5421;
    reg [7:0] z5421_assgn54210;
    reg [7:0] z5421_assgn54211;
    reg [7:0] z5421_assgn54212;
    reg [7:0] z5421_assgn54213;
    reg [7:0] z2035_assgn2035;
    wire [7:0] p3_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5439_assgn5439;
    reg [7:0] z5439_assgn54390;
    reg [7:0] z5439_assgn54391;
    reg [7:0] z5439_assgn54392;
    reg [7:0] z5439_assgn54393;
    reg [7:0] z2051_assgn2051;
    wire [7:0] u0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5443_assgn5443;
    reg [7:0] z5443_assgn54430;
    reg [7:0] z5443_assgn54431;
    reg [7:0] z5443_assgn54432;
    reg [7:0] z5443_assgn54433;
    reg [7:0] z2053_assgn2053;
    wire [7:0] u1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5451_assgn5451;
    reg [7:0] z5451_assgn54510;
    reg [7:0] z5451_assgn54511;
    reg [7:0] z5451_assgn54512;
    reg [7:0] z5451_assgn54513;
    reg [7:0] z2059_assgn2059;
    wire [7:0] p0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5455_assgn5455;
    reg [7:0] z5455_assgn54550;
    reg [7:0] z5455_assgn54551;
    reg [7:0] z5455_assgn54552;
    reg [7:0] z5455_assgn54553;
    reg [7:0] z2061_assgn2061;
    wire [7:0] p1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5463_assgn5463;
    reg [7:0] z5463_assgn54630;
    reg [7:0] z5463_assgn54631;
    reg [7:0] z5463_assgn54632;
    reg [7:0] z5463_assgn54633;
    reg [7:0] z2067_assgn2067;
    wire [7:0] p2_hpc22_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5467_assgn5467;
    reg [7:0] z5467_assgn54670;
    reg [7:0] z5467_assgn54671;
    reg [7:0] z5467_assgn54672;
    reg [7:0] z5467_assgn54673;
    reg [7:0] z2069_assgn2069;
    wire [7:0] p3_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul2_G16_mul1_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5479_assgn5479;
    reg [7:0] z5479_assgn54790;
    reg [7:0] z5479_assgn54791;
    reg [7:0] z5479_assgn54792;
    reg [7:0] z5479_assgn54793;
    reg [7:0] z5479_assgn54794;
    reg [7:0] z2079_assgn2079;
    wire [7:0] p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] z5483_assgn5483;
    reg [7:0] z5483_assgn54830;
    reg [7:0] z5483_assgn54831;
    reg [7:0] z5483_assgn54832;
    reg [7:0] z5483_assgn54833;
    reg [7:0] z5483_assgn54834;
    reg [7:0] z2081_assgn2081;
    wire [7:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G16_mul1_G256_inv0;
    wire [7:0] q0_G16_mul1_G256_inv0;
    wire [7:0] q1_G16_mul1_G256_inv0;
    wire [7:0] z5495_assgn5495;
    reg [7:0] z5495_assgn54950;
    reg [7:0] z5495_assgn54951;
    reg [7:0] z5495_assgn54952;
    reg [7:0] z5495_assgn54953;
    reg [7:0] z5495_assgn54954;
    reg [7:0] z2091_assgn2091;
    wire [7:0] p0ls2_G16_mul1_G256_inv0;
    wire [7:0] z5499_assgn5499;
    reg [7:0] z5499_assgn54990;
    reg [7:0] z5499_assgn54991;
    reg [7:0] z5499_assgn54992;
    reg [7:0] z5499_assgn54993;
    reg [7:0] z5499_assgn54994;
    reg [7:0] z2093_assgn2093;
    wire [7:0] p1ls2_G16_mul1_G256_inv0;
    wire [7:0] p0_G256_inv0;
    wire [7:0] p1_G256_inv0;
    wire [7:0] r00_G16_mul2_G256_inv0;
    wire [7:0] r10_G16_mul2_G256_inv0;
    wire [7:0] r20_G16_mul2_G256_inv0;
    wire [7:0] r30_G16_mul2_G256_inv0;
    wire [7:0] r40_G16_mul2_G256_inv0;
    wire [7:0] r50_G16_mul2_G256_inv0;
    wire [7:0] r60_G16_mul2_G256_inv0;
    wire [7:0] r70_G16_mul2_G256_inv0;
    wire [7:0] r80_G16_mul2_G256_inv0;
    wire [7:0] z5525_assgn5525;
    reg [7:0] z5525_assgn55250;
    reg [7:0] z5525_assgn55251;
    reg [7:0] z5525_assgn55252;
    reg [7:0] z5525_assgn55253;
    reg [7:0] z2117_assgn2117;
    wire [7:0] a0_0_G16_mul2_G256_inv0;
    wire [7:0] z5529_assgn5529;
    reg [7:0] z5529_assgn55290;
    reg [7:0] z5529_assgn55291;
    reg [7:0] z5529_assgn55292;
    reg [7:0] z5529_assgn55293;
    reg [7:0] z2119_assgn2119;
    wire [7:0] a1_0_G16_mul2_G256_inv0;
    wire [7:0] z5533_assgn5533;
    reg [7:0] z5533_assgn55330;
    reg [7:0] z5533_assgn55331;
    reg [7:0] z5533_assgn55332;
    reg [7:0] z5533_assgn55333;
    reg [7:0] z2121_assgn2121;
    wire [7:0] a0_G16_mul2_G256_inv0;
    wire [7:0] z5537_assgn5537;
    reg [7:0] z5537_assgn55370;
    reg [7:0] z5537_assgn55371;
    reg [7:0] z5537_assgn55372;
    reg [7:0] z5537_assgn55373;
    reg [7:0] z2123_assgn2123;
    wire [7:0] a1_G16_mul2_G256_inv0;
    wire [7:0] z5541_assgn5541;
    reg [7:0] z5541_assgn55410;
    reg [7:0] z5541_assgn55411;
    reg [7:0] z5541_assgn55412;
    reg [7:0] z5541_assgn55413;
    reg [7:0] z2125_assgn2125;
    wire [7:0] b0_G16_mul2_G256_inv0;
    wire [7:0] z5545_assgn5545;
    reg [7:0] z5545_assgn55450;
    reg [7:0] z5545_assgn55451;
    reg [7:0] z5545_assgn55452;
    reg [7:0] z5545_assgn55453;
    reg [7:0] z2127_assgn2127;
    wire [7:0] b1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G16_mul2_G256_inv0;
    wire [7:0] c0_G16_mul2_G256_inv0;
    wire [7:0] c1_G16_mul2_G256_inv0;
    wire [7:0] d0_G16_mul2_G256_inv0;
    wire [7:0] d1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5575_assgn5575;
    reg [7:0] z5575_assgn55750;
    reg [7:0] z5575_assgn55751;
    reg [7:0] z5575_assgn55752;
    reg [7:0] z5575_assgn55753;
    reg [7:0] z2155_assgn2155;
    wire [7:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5579_assgn5579;
    reg [7:0] z5579_assgn55790;
    reg [7:0] z5579_assgn55791;
    reg [7:0] z5579_assgn55792;
    reg [7:0] z5579_assgn55793;
    reg [7:0] z2157_assgn2157;
    wire [7:0] a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5583_assgn5583;
    reg [7:0] z5583_assgn55830;
    reg [7:0] z5583_assgn55831;
    reg [7:0] z5583_assgn55832;
    reg [7:0] z5583_assgn55833;
    reg [7:0] z2159_assgn2159;
    wire [7:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5587_assgn5587;
    reg [7:0] z5587_assgn55870;
    reg [7:0] z5587_assgn55871;
    reg [7:0] z5587_assgn55872;
    reg [7:0] z5587_assgn55873;
    reg [7:0] z2161_assgn2161;
    wire [7:0] a1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5591_assgn5591;
    reg [7:0] z5591_assgn55910;
    reg [7:0] z5591_assgn55911;
    reg [7:0] z5591_assgn55912;
    reg [7:0] z5591_assgn55913;
    reg [7:0] z2163_assgn2163;
    wire [7:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5595_assgn5595;
    reg [7:0] z5595_assgn55950;
    reg [7:0] z5595_assgn55951;
    reg [7:0] z5595_assgn55952;
    reg [7:0] z5595_assgn55953;
    reg [7:0] z2165_assgn2165;
    wire [7:0] b1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5625_assgn5625;
    reg [7:0] z5625_assgn56250;
    reg [7:0] z5625_assgn56251;
    reg [7:0] z5625_assgn56252;
    reg [7:0] z5625_assgn56253;
    reg [7:0] z2193_assgn2193;
    wire [7:0] u0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5629_assgn5629;
    reg [7:0] z5629_assgn56290;
    reg [7:0] z5629_assgn56291;
    reg [7:0] z5629_assgn56292;
    reg [7:0] z5629_assgn56293;
    reg [7:0] z2195_assgn2195;
    wire [7:0] u1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5637_assgn5637;
    reg [7:0] z5637_assgn56370;
    reg [7:0] z5637_assgn56371;
    reg [7:0] z5637_assgn56372;
    reg [7:0] z5637_assgn56373;
    reg [7:0] z2201_assgn2201;
    wire [7:0] p0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5641_assgn5641;
    reg [7:0] z5641_assgn56410;
    reg [7:0] z5641_assgn56411;
    reg [7:0] z5641_assgn56412;
    reg [7:0] z5641_assgn56413;
    reg [7:0] z2203_assgn2203;
    wire [7:0] p1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5649_assgn5649;
    reg [7:0] z5649_assgn56490;
    reg [7:0] z5649_assgn56491;
    reg [7:0] z5649_assgn56492;
    reg [7:0] z5649_assgn56493;
    reg [7:0] z2209_assgn2209;
    wire [7:0] p2_hpc20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5653_assgn5653;
    reg [7:0] z5653_assgn56530;
    reg [7:0] z5653_assgn56531;
    reg [7:0] z5653_assgn56532;
    reg [7:0] z5653_assgn56533;
    reg [7:0] z2211_assgn2211;
    wire [7:0] p3_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5667_assgn5667;
    reg [7:0] z5667_assgn56670;
    reg [7:0] z5667_assgn56671;
    reg [7:0] z5667_assgn56672;
    reg [7:0] z5667_assgn56673;
    reg [7:0] z2223_assgn2223;
    wire [7:0] u0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5671_assgn5671;
    reg [7:0] z5671_assgn56710;
    reg [7:0] z5671_assgn56711;
    reg [7:0] z5671_assgn56712;
    reg [7:0] z5671_assgn56713;
    reg [7:0] z2225_assgn2225;
    wire [7:0] u1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5679_assgn5679;
    reg [7:0] z5679_assgn56790;
    reg [7:0] z5679_assgn56791;
    reg [7:0] z5679_assgn56792;
    reg [7:0] z5679_assgn56793;
    reg [7:0] z2231_assgn2231;
    wire [7:0] p0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5683_assgn5683;
    reg [7:0] z5683_assgn56830;
    reg [7:0] z5683_assgn56831;
    reg [7:0] z5683_assgn56832;
    reg [7:0] z5683_assgn56833;
    reg [7:0] z2233_assgn2233;
    wire [7:0] p1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5691_assgn5691;
    reg [7:0] z5691_assgn56910;
    reg [7:0] z5691_assgn56911;
    reg [7:0] z5691_assgn56912;
    reg [7:0] z5691_assgn56913;
    reg [7:0] z2239_assgn2239;
    wire [7:0] p2_hpc21_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5695_assgn5695;
    reg [7:0] z5695_assgn56950;
    reg [7:0] z5695_assgn56951;
    reg [7:0] z5695_assgn56952;
    reg [7:0] z5695_assgn56953;
    reg [7:0] z2241_assgn2241;
    wire [7:0] p3_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5713_assgn5713;
    reg [7:0] z5713_assgn57130;
    reg [7:0] z5713_assgn57131;
    reg [7:0] z5713_assgn57132;
    reg [7:0] z5713_assgn57133;
    reg [7:0] z2257_assgn2257;
    wire [7:0] u0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5717_assgn5717;
    reg [7:0] z5717_assgn57170;
    reg [7:0] z5717_assgn57171;
    reg [7:0] z5717_assgn57172;
    reg [7:0] z5717_assgn57173;
    reg [7:0] z2259_assgn2259;
    wire [7:0] u1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5725_assgn5725;
    reg [7:0] z5725_assgn57250;
    reg [7:0] z5725_assgn57251;
    reg [7:0] z5725_assgn57252;
    reg [7:0] z5725_assgn57253;
    reg [7:0] z2265_assgn2265;
    wire [7:0] p0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5729_assgn5729;
    reg [7:0] z5729_assgn57290;
    reg [7:0] z5729_assgn57291;
    reg [7:0] z5729_assgn57292;
    reg [7:0] z5729_assgn57293;
    reg [7:0] z2267_assgn2267;
    wire [7:0] p1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5737_assgn5737;
    reg [7:0] z5737_assgn57370;
    reg [7:0] z5737_assgn57371;
    reg [7:0] z5737_assgn57372;
    reg [7:0] z5737_assgn57373;
    reg [7:0] z2273_assgn2273;
    wire [7:0] p2_hpc22_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5741_assgn5741;
    reg [7:0] z5741_assgn57410;
    reg [7:0] z5741_assgn57411;
    reg [7:0] z5741_assgn57412;
    reg [7:0] z5741_assgn57413;
    reg [7:0] z2275_assgn2275;
    wire [7:0] p3_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul0_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5753_assgn5753;
    reg [7:0] z5753_assgn57530;
    reg [7:0] z5753_assgn57531;
    reg [7:0] z5753_assgn57532;
    reg [7:0] z5753_assgn57533;
    reg [7:0] z5753_assgn57534;
    reg [7:0] z2285_assgn2285;
    wire [7:0] p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] z5757_assgn5757;
    reg [7:0] z5757_assgn57570;
    reg [7:0] z5757_assgn57571;
    reg [7:0] z5757_assgn57572;
    reg [7:0] z5757_assgn57573;
    reg [7:0] z5757_assgn57574;
    reg [7:0] z2287_assgn2287;
    wire [7:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G16_mul2_G256_inv0;
    wire [7:0] e1_G16_mul2_G256_inv0;
    wire [7:0] z5765_assgn5765;
    reg [7:0] z5765_assgn57650;
    reg [7:0] z5765_assgn57651;
    reg [7:0] z5765_assgn57652;
    reg [7:0] z5765_assgn57653;
    reg [7:0] z5765_assgn57654;
    reg [7:0] z2293_assgn2293;
    wire [7:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5769_assgn5769;
    reg [7:0] z5769_assgn57690;
    reg [7:0] z5769_assgn57691;
    reg [7:0] z5769_assgn57692;
    reg [7:0] z5769_assgn57693;
    reg [7:0] z5769_assgn57694;
    reg [7:0] z2295_assgn2295;
    wire [7:0] a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5773_assgn5773;
    reg [7:0] z5773_assgn57730;
    reg [7:0] z5773_assgn57731;
    reg [7:0] z5773_assgn57732;
    reg [7:0] z5773_assgn57733;
    reg [7:0] z5773_assgn57734;
    reg [7:0] z2297_assgn2297;
    wire [7:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5777_assgn5777;
    reg [7:0] z5777_assgn57770;
    reg [7:0] z5777_assgn57771;
    reg [7:0] z5777_assgn57772;
    reg [7:0] z5777_assgn57773;
    reg [7:0] z5777_assgn57774;
    reg [7:0] z2299_assgn2299;
    wire [7:0] a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5781_assgn5781;
    reg [7:0] z5781_assgn57810;
    reg [7:0] z5781_assgn57811;
    reg [7:0] z5781_assgn57812;
    reg [7:0] z5781_assgn57813;
    reg [7:0] z5781_assgn57814;
    reg [7:0] z2301_assgn2301;
    wire [7:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5785_assgn5785;
    reg [7:0] z5785_assgn57850;
    reg [7:0] z5785_assgn57851;
    reg [7:0] z5785_assgn57852;
    reg [7:0] z5785_assgn57853;
    reg [7:0] z5785_assgn57854;
    reg [7:0] z2303_assgn2303;
    wire [7:0] b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5797_assgn5797;
    reg [7:0] z5797_assgn57970;
    reg [7:0] z5797_assgn57971;
    reg [7:0] z5797_assgn57972;
    reg [7:0] z5797_assgn57973;
    reg [7:0] z5797_assgn57974;
    reg [7:0] z2313_assgn2313;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] z5801_assgn5801;
    reg [7:0] z5801_assgn58010;
    reg [7:0] z5801_assgn58011;
    reg [7:0] z5801_assgn58012;
    reg [7:0] z5801_assgn58013;
    reg [7:0] z5801_assgn58014;
    reg [7:0] z2315_assgn2315;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] e01_G16_mul2_G256_inv0;
    wire [7:0] e11_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5815_assgn5815;
    reg [7:0] z5815_assgn58150;
    reg [7:0] z5815_assgn58151;
    reg [7:0] z5815_assgn58152;
    reg [7:0] z5815_assgn58153;
    reg [7:0] z2327_assgn2327;
    wire [7:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5819_assgn5819;
    reg [7:0] z5819_assgn58190;
    reg [7:0] z5819_assgn58191;
    reg [7:0] z5819_assgn58192;
    reg [7:0] z5819_assgn58193;
    reg [7:0] z2329_assgn2329;
    wire [7:0] a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5823_assgn5823;
    reg [7:0] z5823_assgn58230;
    reg [7:0] z5823_assgn58231;
    reg [7:0] z5823_assgn58232;
    reg [7:0] z5823_assgn58233;
    reg [7:0] z2331_assgn2331;
    wire [7:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5827_assgn5827;
    reg [7:0] z5827_assgn58270;
    reg [7:0] z5827_assgn58271;
    reg [7:0] z5827_assgn58272;
    reg [7:0] z5827_assgn58273;
    reg [7:0] z2333_assgn2333;
    wire [7:0] a1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5831_assgn5831;
    reg [7:0] z5831_assgn58310;
    reg [7:0] z5831_assgn58311;
    reg [7:0] z5831_assgn58312;
    reg [7:0] z5831_assgn58313;
    reg [7:0] z2335_assgn2335;
    wire [7:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5835_assgn5835;
    reg [7:0] z5835_assgn58350;
    reg [7:0] z5835_assgn58351;
    reg [7:0] z5835_assgn58352;
    reg [7:0] z5835_assgn58353;
    reg [7:0] z2337_assgn2337;
    wire [7:0] b1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5865_assgn5865;
    reg [7:0] z5865_assgn58650;
    reg [7:0] z5865_assgn58651;
    reg [7:0] z5865_assgn58652;
    reg [7:0] z5865_assgn58653;
    reg [7:0] z2365_assgn2365;
    wire [7:0] u0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5869_assgn5869;
    reg [7:0] z5869_assgn58690;
    reg [7:0] z5869_assgn58691;
    reg [7:0] z5869_assgn58692;
    reg [7:0] z5869_assgn58693;
    reg [7:0] z2367_assgn2367;
    wire [7:0] u1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5877_assgn5877;
    reg [7:0] z5877_assgn58770;
    reg [7:0] z5877_assgn58771;
    reg [7:0] z5877_assgn58772;
    reg [7:0] z5877_assgn58773;
    reg [7:0] z2373_assgn2373;
    wire [7:0] p0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5881_assgn5881;
    reg [7:0] z5881_assgn58810;
    reg [7:0] z5881_assgn58811;
    reg [7:0] z5881_assgn58812;
    reg [7:0] z5881_assgn58813;
    reg [7:0] z2375_assgn2375;
    wire [7:0] p1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5889_assgn5889;
    reg [7:0] z5889_assgn58890;
    reg [7:0] z5889_assgn58891;
    reg [7:0] z5889_assgn58892;
    reg [7:0] z5889_assgn58893;
    reg [7:0] z2381_assgn2381;
    wire [7:0] p2_hpc20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5893_assgn5893;
    reg [7:0] z5893_assgn58930;
    reg [7:0] z5893_assgn58931;
    reg [7:0] z5893_assgn58932;
    reg [7:0] z5893_assgn58933;
    reg [7:0] z2383_assgn2383;
    wire [7:0] p3_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5907_assgn5907;
    reg [7:0] z5907_assgn59070;
    reg [7:0] z5907_assgn59071;
    reg [7:0] z5907_assgn59072;
    reg [7:0] z5907_assgn59073;
    reg [7:0] z2395_assgn2395;
    wire [7:0] u0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5911_assgn5911;
    reg [7:0] z5911_assgn59110;
    reg [7:0] z5911_assgn59111;
    reg [7:0] z5911_assgn59112;
    reg [7:0] z5911_assgn59113;
    reg [7:0] z2397_assgn2397;
    wire [7:0] u1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5919_assgn5919;
    reg [7:0] z5919_assgn59190;
    reg [7:0] z5919_assgn59191;
    reg [7:0] z5919_assgn59192;
    reg [7:0] z5919_assgn59193;
    reg [7:0] z2403_assgn2403;
    wire [7:0] p0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5923_assgn5923;
    reg [7:0] z5923_assgn59230;
    reg [7:0] z5923_assgn59231;
    reg [7:0] z5923_assgn59232;
    reg [7:0] z5923_assgn59233;
    reg [7:0] z2405_assgn2405;
    wire [7:0] p1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5931_assgn5931;
    reg [7:0] z5931_assgn59310;
    reg [7:0] z5931_assgn59311;
    reg [7:0] z5931_assgn59312;
    reg [7:0] z5931_assgn59313;
    reg [7:0] z2411_assgn2411;
    wire [7:0] p2_hpc21_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5935_assgn5935;
    reg [7:0] z5935_assgn59350;
    reg [7:0] z5935_assgn59351;
    reg [7:0] z5935_assgn59352;
    reg [7:0] z5935_assgn59353;
    reg [7:0] z2413_assgn2413;
    wire [7:0] p3_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5953_assgn5953;
    reg [7:0] z5953_assgn59530;
    reg [7:0] z5953_assgn59531;
    reg [7:0] z5953_assgn59532;
    reg [7:0] z5953_assgn59533;
    reg [7:0] z2429_assgn2429;
    wire [7:0] u0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5957_assgn5957;
    reg [7:0] z5957_assgn59570;
    reg [7:0] z5957_assgn59571;
    reg [7:0] z5957_assgn59572;
    reg [7:0] z5957_assgn59573;
    reg [7:0] z2431_assgn2431;
    wire [7:0] u1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5965_assgn5965;
    reg [7:0] z5965_assgn59650;
    reg [7:0] z5965_assgn59651;
    reg [7:0] z5965_assgn59652;
    reg [7:0] z5965_assgn59653;
    reg [7:0] z2437_assgn2437;
    wire [7:0] p0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5969_assgn5969;
    reg [7:0] z5969_assgn59690;
    reg [7:0] z5969_assgn59691;
    reg [7:0] z5969_assgn59692;
    reg [7:0] z5969_assgn59693;
    reg [7:0] z2439_assgn2439;
    wire [7:0] p1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5977_assgn5977;
    reg [7:0] z5977_assgn59770;
    reg [7:0] z5977_assgn59771;
    reg [7:0] z5977_assgn59772;
    reg [7:0] z5977_assgn59773;
    reg [7:0] z2445_assgn2445;
    wire [7:0] p2_hpc22_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5981_assgn5981;
    reg [7:0] z5981_assgn59810;
    reg [7:0] z5981_assgn59811;
    reg [7:0] z5981_assgn59812;
    reg [7:0] z5981_assgn59813;
    reg [7:0] z2447_assgn2447;
    wire [7:0] p3_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul1_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5993_assgn5993;
    reg [7:0] z5993_assgn59930;
    reg [7:0] z5993_assgn59931;
    reg [7:0] z5993_assgn59932;
    reg [7:0] z5993_assgn59933;
    reg [7:0] z5993_assgn59934;
    reg [7:0] z2457_assgn2457;
    wire [7:0] p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] z5997_assgn5997;
    reg [7:0] z5997_assgn59970;
    reg [7:0] z5997_assgn59971;
    reg [7:0] z5997_assgn59972;
    reg [7:0] z5997_assgn59973;
    reg [7:0] z5997_assgn59974;
    reg [7:0] z2459_assgn2459;
    wire [7:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G16_mul2_G256_inv0;
    wire [7:0] p0_G16_mul2_G256_inv0;
    wire [7:0] p1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6015_assgn6015;
    reg [7:0] z6015_assgn60150;
    reg [7:0] z6015_assgn60151;
    reg [7:0] z6015_assgn60152;
    reg [7:0] z6015_assgn60153;
    reg [7:0] z2475_assgn2475;
    wire [7:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6019_assgn6019;
    reg [7:0] z6019_assgn60190;
    reg [7:0] z6019_assgn60191;
    reg [7:0] z6019_assgn60192;
    reg [7:0] z6019_assgn60193;
    reg [7:0] z2477_assgn2477;
    wire [7:0] a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6023_assgn6023;
    reg [7:0] z6023_assgn60230;
    reg [7:0] z6023_assgn60231;
    reg [7:0] z6023_assgn60232;
    reg [7:0] z6023_assgn60233;
    reg [7:0] z2479_assgn2479;
    wire [7:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6027_assgn6027;
    reg [7:0] z6027_assgn60270;
    reg [7:0] z6027_assgn60271;
    reg [7:0] z6027_assgn60272;
    reg [7:0] z6027_assgn60273;
    reg [7:0] z2481_assgn2481;
    wire [7:0] a1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6031_assgn6031;
    reg [7:0] z6031_assgn60310;
    reg [7:0] z6031_assgn60311;
    reg [7:0] z6031_assgn60312;
    reg [7:0] z6031_assgn60313;
    reg [7:0] z2483_assgn2483;
    wire [7:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6035_assgn6035;
    reg [7:0] z6035_assgn60350;
    reg [7:0] z6035_assgn60351;
    reg [7:0] z6035_assgn60352;
    reg [7:0] z6035_assgn60353;
    reg [7:0] z2485_assgn2485;
    wire [7:0] b1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6065_assgn6065;
    reg [7:0] z6065_assgn60650;
    reg [7:0] z6065_assgn60651;
    reg [7:0] z6065_assgn60652;
    reg [7:0] z6065_assgn60653;
    reg [7:0] z2513_assgn2513;
    wire [7:0] u0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6069_assgn6069;
    reg [7:0] z6069_assgn60690;
    reg [7:0] z6069_assgn60691;
    reg [7:0] z6069_assgn60692;
    reg [7:0] z6069_assgn60693;
    reg [7:0] z2515_assgn2515;
    wire [7:0] u1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6077_assgn6077;
    reg [7:0] z6077_assgn60770;
    reg [7:0] z6077_assgn60771;
    reg [7:0] z6077_assgn60772;
    reg [7:0] z6077_assgn60773;
    reg [7:0] z2521_assgn2521;
    wire [7:0] p0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6081_assgn6081;
    reg [7:0] z6081_assgn60810;
    reg [7:0] z6081_assgn60811;
    reg [7:0] z6081_assgn60812;
    reg [7:0] z6081_assgn60813;
    reg [7:0] z2523_assgn2523;
    wire [7:0] p1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] e0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6089_assgn6089;
    reg [7:0] z6089_assgn60890;
    reg [7:0] z6089_assgn60891;
    reg [7:0] z6089_assgn60892;
    reg [7:0] z6089_assgn60893;
    reg [7:0] z2529_assgn2529;
    wire [7:0] p2_hpc20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6093_assgn6093;
    reg [7:0] z6093_assgn60930;
    reg [7:0] z6093_assgn60931;
    reg [7:0] z6093_assgn60932;
    reg [7:0] z6093_assgn60933;
    reg [7:0] z2531_assgn2531;
    wire [7:0] p3_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc20_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] e1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6107_assgn6107;
    reg [7:0] z6107_assgn61070;
    reg [7:0] z6107_assgn61071;
    reg [7:0] z6107_assgn61072;
    reg [7:0] z6107_assgn61073;
    reg [7:0] z2543_assgn2543;
    wire [7:0] u0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6111_assgn6111;
    reg [7:0] z6111_assgn61110;
    reg [7:0] z6111_assgn61111;
    reg [7:0] z6111_assgn61112;
    reg [7:0] z6111_assgn61113;
    reg [7:0] z2545_assgn2545;
    wire [7:0] u1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6119_assgn6119;
    reg [7:0] z6119_assgn61190;
    reg [7:0] z6119_assgn61191;
    reg [7:0] z6119_assgn61192;
    reg [7:0] z6119_assgn61193;
    reg [7:0] z2551_assgn2551;
    wire [7:0] p0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6123_assgn6123;
    reg [7:0] z6123_assgn61230;
    reg [7:0] z6123_assgn61231;
    reg [7:0] z6123_assgn61232;
    reg [7:0] z6123_assgn61233;
    reg [7:0] z2553_assgn2553;
    wire [7:0] p1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6131_assgn6131;
    reg [7:0] z6131_assgn61310;
    reg [7:0] z6131_assgn61311;
    reg [7:0] z6131_assgn61312;
    reg [7:0] z6131_assgn61313;
    reg [7:0] z2559_assgn2559;
    wire [7:0] p2_hpc21_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6135_assgn6135;
    reg [7:0] z6135_assgn61350;
    reg [7:0] z6135_assgn61351;
    reg [7:0] z6135_assgn61352;
    reg [7:0] z6135_assgn61353;
    reg [7:0] z2561_assgn2561;
    wire [7:0] p3_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc21_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6153_assgn6153;
    reg [7:0] z6153_assgn61530;
    reg [7:0] z6153_assgn61531;
    reg [7:0] z6153_assgn61532;
    reg [7:0] z6153_assgn61533;
    reg [7:0] z2577_assgn2577;
    wire [7:0] u0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6157_assgn6157;
    reg [7:0] z6157_assgn61570;
    reg [7:0] z6157_assgn61571;
    reg [7:0] z6157_assgn61572;
    reg [7:0] z6157_assgn61573;
    reg [7:0] z2579_assgn2579;
    wire [7:0] u1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] v1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6165_assgn6165;
    reg [7:0] z6165_assgn61650;
    reg [7:0] z6165_assgn61651;
    reg [7:0] z6165_assgn61652;
    reg [7:0] z6165_assgn61653;
    reg [7:0] z2585_assgn2585;
    wire [7:0] p0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6169_assgn6169;
    reg [7:0] z6169_assgn61690;
    reg [7:0] z6169_assgn61691;
    reg [7:0] z6169_assgn61692;
    reg [7:0] z6169_assgn61693;
    reg [7:0] z2587_assgn2587;
    wire [7:0] p1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p01_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6177_assgn6177;
    reg [7:0] z6177_assgn61770;
    reg [7:0] z6177_assgn61771;
    reg [7:0] z6177_assgn61772;
    reg [7:0] z6177_assgn61773;
    reg [7:0] z2593_assgn2593;
    wire [7:0] p2_hpc22_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6181_assgn6181;
    reg [7:0] z6181_assgn61810;
    reg [7:0] z6181_assgn61811;
    reg [7:0] z6181_assgn61812;
    reg [7:0] z6181_assgn61813;
    reg [7:0] z2595_assgn2595;
    wire [7:0] p3_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [7:0] p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] p23_hpc22_G4_mul2_G16_mul2_G256_inv0;
    reg [7:0] p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [7:0] q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6193_assgn6193;
    reg [7:0] z6193_assgn61930;
    reg [7:0] z6193_assgn61931;
    reg [7:0] z6193_assgn61932;
    reg [7:0] z6193_assgn61933;
    reg [7:0] z6193_assgn61934;
    reg [7:0] z2605_assgn2605;
    wire [7:0] p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] z6197_assgn6197;
    reg [7:0] z6197_assgn61970;
    reg [7:0] z6197_assgn61971;
    reg [7:0] z6197_assgn61972;
    reg [7:0] z6197_assgn61973;
    reg [7:0] z6197_assgn61974;
    reg [7:0] z2607_assgn2607;
    wire [7:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G16_mul2_G256_inv0;
    wire [7:0] q0_G16_mul2_G256_inv0;
    wire [7:0] q1_G16_mul2_G256_inv0;
    wire [7:0] z6209_assgn6209;
    reg [7:0] z6209_assgn62090;
    reg [7:0] z6209_assgn62091;
    reg [7:0] z6209_assgn62092;
    reg [7:0] z6209_assgn62093;
    reg [7:0] z6209_assgn62094;
    reg [7:0] z2617_assgn2617;
    wire [7:0] p0ls2_G16_mul2_G256_inv0;
    wire [7:0] z6213_assgn6213;
    reg [7:0] z6213_assgn62130;
    reg [7:0] z6213_assgn62131;
    reg [7:0] z6213_assgn62132;
    reg [7:0] z6213_assgn62133;
    reg [7:0] z6213_assgn62134;
    reg [7:0] z2619_assgn2619;
    wire [7:0] p1ls2_G16_mul2_G256_inv0;
    wire [7:0] q0_G256_inv0;
    wire [7:0] q1_G256_inv0;
    wire [7:0] z6221_assgn6221;
    reg [7:0] z6221_assgn62210;
    reg [7:0] z6221_assgn62211;
    reg [7:0] z6221_assgn62212;
    reg [7:0] z6221_assgn62213;
    reg [7:0] z6221_assgn62214;
    reg [7:0] z2625_assgn2625;
    wire [7:0] p0ls4_G256_inv0;
    wire [7:0] z6225_assgn6225;
    reg [7:0] z6225_assgn62250;
    reg [7:0] z6225_assgn62251;
    reg [7:0] z6225_assgn62252;
    reg [7:0] z6225_assgn62253;
    reg [7:0] z6225_assgn62254;
    reg [7:0] z2627_assgn2627;
    wire [7:0] p1ls4_G256_inv0;
    wire [7:0] t4;
    wire [7:0] t5;
    wire [7:0] y_G256_newbasis1;
    wire [7:0] tempy1_G256_newbasis1;
    wire [7:0] z6237_assgn6237;
    reg [7:0] z6237_assgn62370;
    reg [7:0] z6237_assgn62371;
    reg [7:0] z6237_assgn62372;
    reg [7:0] z6237_assgn62373;
    reg [7:0] z6237_assgn62374;
    reg [7:0] z2637_assgn2637;
    wire [7:0] cond1_G256_newbasis1;
    wire [7:0] negCond1_G256_newbasis1;
    wire [7:0] yxorb1_G256_newbasis1;
    wire [7:0] z6245_assgn6245;
    reg [7:0] z6245_assgn62450;
    reg [7:0] z6245_assgn62451;
    reg [7:0] z6245_assgn62452;
    reg [7:0] z6245_assgn62453;
    reg [7:0] z6245_assgn62454;
    reg [7:0] z2643_assgn2643;
    wire [7:0] ny1_G256_newbasis1;
    wire [7:0] z6249_assgn6249;
    reg [7:0] z6249_assgn62490;
    reg [7:0] z6249_assgn62491;
    reg [7:0] z6249_assgn62492;
    reg [7:0] z6249_assgn62493;
    reg [7:0] z6249_assgn62494;
    reg [7:0] z2646_assgn2646;
    wire [7:0] tempyIntoNegCond1_G256_newbasis1;
    wire [7:0] y1_G256_newbasis1;
    wire [7:0] z6255_assgn6255;
    reg [7:0] z6255_assgn62550;
    reg [7:0] z6255_assgn62551;
    reg [7:0] z6255_assgn62552;
    reg [7:0] z6255_assgn62553;
    reg [7:0] z6255_assgn62554;
    reg [7:0] z2649_assgn2649;
    wire [7:0] x1_G256_newbasis1;
    wire [7:0] tempy2_G256_newbasis1;
    wire [7:0] z6261_assgn6261;
    reg [7:0] z6261_assgn62610;
    reg [7:0] z6261_assgn62611;
    reg [7:0] z6261_assgn62612;
    reg [7:0] z6261_assgn62613;
    reg [7:0] z6261_assgn62614;
    reg [7:0] z2653_assgn2653;
    wire [7:0] cond2_G256_newbasis1;
    wire [7:0] negCond2_G256_newbasis1;
    wire [7:0] z6267_assgn6267;
    reg [7:0] z6267_assgn62670;
    reg [7:0] z6267_assgn62671;
    reg [7:0] z6267_assgn62672;
    reg [7:0] z6267_assgn62673;
    reg [7:0] z6267_assgn62674;
    reg [7:0] z2657_assgn2657;
    wire [7:0] yxorb2_G256_newbasis1;
    wire [7:0] ny2_G256_newbasis1;
    wire [7:0] tempyIntoNegCond2_G256_newbasis1;
    wire [7:0] y2_G256_newbasis1;
    wire [7:0] z6277_assgn6277;
    reg [7:0] z6277_assgn62770;
    reg [7:0] z6277_assgn62771;
    reg [7:0] z6277_assgn62772;
    reg [7:0] z6277_assgn62773;
    reg [7:0] z6277_assgn62774;
    reg [7:0] z2665_assgn2665;
    wire [7:0] x2_G256_newbasis1;
    wire [7:0] tempy3_G256_newbasis1;
    wire [7:0] z6283_assgn6283;
    reg [7:0] z6283_assgn62830;
    reg [7:0] z6283_assgn62831;
    reg [7:0] z6283_assgn62832;
    reg [7:0] z6283_assgn62833;
    reg [7:0] z6283_assgn62834;
    reg [7:0] z2669_assgn2669;
    wire [7:0] cond3_G256_newbasis1;
    wire [7:0] negCond3_G256_newbasis1;
    wire [7:0] z6289_assgn6289;
    reg [7:0] z6289_assgn62890;
    reg [7:0] z6289_assgn62891;
    reg [7:0] z6289_assgn62892;
    reg [7:0] z6289_assgn62893;
    reg [7:0] z6289_assgn62894;
    reg [7:0] z2673_assgn2673;
    wire [7:0] yxorb3_G256_newbasis1;
    wire [7:0] ny3_G256_newbasis1;
    wire [7:0] tempyIntoNegCond3_G256_newbasis1;
    wire [7:0] y3_G256_newbasis1;
    wire [7:0] z6299_assgn6299;
    reg [7:0] z6299_assgn62990;
    reg [7:0] z6299_assgn62991;
    reg [7:0] z6299_assgn62992;
    reg [7:0] z6299_assgn62993;
    reg [7:0] z6299_assgn62994;
    reg [7:0] z2681_assgn2681;
    wire [7:0] x3_G256_newbasis1;
    wire [7:0] tempy4_G256_newbasis1;
    wire [7:0] z6305_assgn6305;
    reg [7:0] z6305_assgn63050;
    reg [7:0] z6305_assgn63051;
    reg [7:0] z6305_assgn63052;
    reg [7:0] z6305_assgn63053;
    reg [7:0] z6305_assgn63054;
    reg [7:0] z2685_assgn2685;
    wire [7:0] cond4_G256_newbasis1;
    wire [7:0] negCond4_G256_newbasis1;
    wire [7:0] z6311_assgn6311;
    reg [7:0] z6311_assgn63110;
    reg [7:0] z6311_assgn63111;
    reg [7:0] z6311_assgn63112;
    reg [7:0] z6311_assgn63113;
    reg [7:0] z6311_assgn63114;
    reg [7:0] z2689_assgn2689;
    wire [7:0] yxorb4_G256_newbasis1;
    wire [7:0] ny4_G256_newbasis1;
    wire [7:0] tempyIntoNegCond4_G256_newbasis1;
    wire [7:0] y4_G256_newbasis1;
    wire [7:0] z6321_assgn6321;
    reg [7:0] z6321_assgn63210;
    reg [7:0] z6321_assgn63211;
    reg [7:0] z6321_assgn63212;
    reg [7:0] z6321_assgn63213;
    reg [7:0] z6321_assgn63214;
    reg [7:0] z2697_assgn2697;
    wire [7:0] x4_G256_newbasis1;
    wire [7:0] tempy5_G256_newbasis1;
    wire [7:0] z6327_assgn6327;
    reg [7:0] z6327_assgn63270;
    reg [7:0] z6327_assgn63271;
    reg [7:0] z6327_assgn63272;
    reg [7:0] z6327_assgn63273;
    reg [7:0] z6327_assgn63274;
    reg [7:0] z2701_assgn2701;
    wire [7:0] cond5_G256_newbasis1;
    wire [7:0] negCond5_G256_newbasis1;
    wire [7:0] z6333_assgn6333;
    reg [7:0] z6333_assgn63330;
    reg [7:0] z6333_assgn63331;
    reg [7:0] z6333_assgn63332;
    reg [7:0] z6333_assgn63333;
    reg [7:0] z6333_assgn63334;
    reg [7:0] z2705_assgn2705;
    wire [7:0] yxorb5_G256_newbasis1;
    wire [7:0] ny5_G256_newbasis1;
    wire [7:0] tempyIntoNegCond5_G256_newbasis1;
    wire [7:0] y5_G256_newbasis1;
    wire [7:0] z6343_assgn6343;
    reg [7:0] z6343_assgn63430;
    reg [7:0] z6343_assgn63431;
    reg [7:0] z6343_assgn63432;
    reg [7:0] z6343_assgn63433;
    reg [7:0] z6343_assgn63434;
    reg [7:0] z2713_assgn2713;
    wire [7:0] x5_G256_newbasis1;
    wire [7:0] tempy6_G256_newbasis1;
    wire [7:0] z6349_assgn6349;
    reg [7:0] z6349_assgn63490;
    reg [7:0] z6349_assgn63491;
    reg [7:0] z6349_assgn63492;
    reg [7:0] z6349_assgn63493;
    reg [7:0] z6349_assgn63494;
    reg [7:0] z2717_assgn2717;
    wire [7:0] cond6_G256_newbasis1;
    wire [7:0] negCond6_G256_newbasis1;
    wire [7:0] z6355_assgn6355;
    reg [7:0] z6355_assgn63550;
    reg [7:0] z6355_assgn63551;
    reg [7:0] z6355_assgn63552;
    reg [7:0] z6355_assgn63553;
    reg [7:0] z6355_assgn63554;
    reg [7:0] z2721_assgn2721;
    wire [7:0] yxorb6_G256_newbasis1;
    wire [7:0] ny6_G256_newbasis1;
    wire [7:0] tempyIntoNegCond6_G256_newbasis1;
    wire [7:0] y6_G256_newbasis1;
    wire [7:0] z6365_assgn6365;
    reg [7:0] z6365_assgn63650;
    reg [7:0] z6365_assgn63651;
    reg [7:0] z6365_assgn63652;
    reg [7:0] z6365_assgn63653;
    reg [7:0] z6365_assgn63654;
    reg [7:0] z2729_assgn2729;
    wire [7:0] x6_G256_newbasis1;
    wire [7:0] tempy7_G256_newbasis1;
    wire [7:0] z6371_assgn6371;
    reg [7:0] z6371_assgn63710;
    reg [7:0] z6371_assgn63711;
    reg [7:0] z6371_assgn63712;
    reg [7:0] z6371_assgn63713;
    reg [7:0] z6371_assgn63714;
    reg [7:0] z2733_assgn2733;
    wire [7:0] cond7_G256_newbasis1;
    wire [7:0] negCond7_G256_newbasis1;
    wire [7:0] z6377_assgn6377;
    reg [7:0] z6377_assgn63770;
    reg [7:0] z6377_assgn63771;
    reg [7:0] z6377_assgn63772;
    reg [7:0] z6377_assgn63773;
    reg [7:0] z6377_assgn63774;
    reg [7:0] z2737_assgn2737;
    wire [7:0] yxorb7_G256_newbasis1;
    wire [7:0] ny7_G256_newbasis1;
    wire [7:0] tempyIntoNegCond7_G256_newbasis1;
    wire [7:0] y7_G256_newbasis1;
    wire [7:0] z6387_assgn6387;
    reg [7:0] z6387_assgn63870;
    reg [7:0] z6387_assgn63871;
    reg [7:0] z6387_assgn63872;
    reg [7:0] z6387_assgn63873;
    reg [7:0] z6387_assgn63874;
    reg [7:0] z2745_assgn2745;
    wire [7:0] x7_G256_newbasis1;
    wire [7:0] tempy8_G256_newbasis1;
    wire [7:0] z6393_assgn6393;
    reg [7:0] z6393_assgn63930;
    reg [7:0] z6393_assgn63931;
    reg [7:0] z6393_assgn63932;
    reg [7:0] z6393_assgn63933;
    reg [7:0] z6393_assgn63934;
    reg [7:0] z2749_assgn2749;
    wire [7:0] cond8_G256_newbasis1;
    wire [7:0] negCond8_G256_newbasis1;
    wire [7:0] z6399_assgn6399;
    reg [7:0] z6399_assgn63990;
    reg [7:0] z6399_assgn63991;
    reg [7:0] z6399_assgn63992;
    reg [7:0] z6399_assgn63993;
    reg [7:0] z6399_assgn63994;
    reg [7:0] z2753_assgn2753;
    wire [7:0] yxorb8_G256_newbasis1;
    wire [7:0] ny8_G256_newbasis1;
    wire [7:0] tempyIntoNegCond8_G256_newbasis1;
    wire [7:0] y8_G256_newbasis1;
    wire [7:0] z6409_assgn6409;
    reg [7:0] z6409_assgn64090;
    reg [7:0] z6409_assgn64091;
    reg [7:0] z6409_assgn64092;
    reg [7:0] z6409_assgn64093;
    reg [7:0] z6409_assgn64094;
    reg [7:0] z2761_assgn2761;
    wire [7:0] x8_G256_newbasis1;
    wire [7:0] t6;
    wire [7:0] z_y_G256_newbasis1;
    wire [7:0] z_tempy1_G256_newbasis1;
    wire [7:0] z6419_assgn6419;
    reg [7:0] z6419_assgn64190;
    reg [7:0] z6419_assgn64191;
    reg [7:0] z6419_assgn64192;
    reg [7:0] z6419_assgn64193;
    reg [7:0] z6419_assgn64194;
    reg [7:0] z2769_assgn2769;
    wire [7:0] z_cond1_G256_newbasis1;
    wire [7:0] z_negCond1_G256_newbasis1;
    wire [7:0] z_yxorb1_G256_newbasis1;
    wire [7:0] z6427_assgn6427;
    reg [7:0] z6427_assgn64270;
    reg [7:0] z6427_assgn64271;
    reg [7:0] z6427_assgn64272;
    reg [7:0] z6427_assgn64273;
    reg [7:0] z6427_assgn64274;
    reg [7:0] z2775_assgn2775;
    wire [7:0] z_ny1_G256_newbasis1;
    wire [7:0] z6431_assgn6431;
    reg [7:0] z6431_assgn64310;
    reg [7:0] z6431_assgn64311;
    reg [7:0] z6431_assgn64312;
    reg [7:0] z6431_assgn64313;
    reg [7:0] z6431_assgn64314;
    reg [7:0] z2778_assgn2778;
    wire [7:0] z_tempyIntoNegCond1_G256_newbasis1;
    wire [7:0] z_y1_G256_newbasis1;
    wire [7:0] z6437_assgn6437;
    reg [7:0] z6437_assgn64370;
    reg [7:0] z6437_assgn64371;
    reg [7:0] z6437_assgn64372;
    reg [7:0] z6437_assgn64373;
    reg [7:0] z6437_assgn64374;
    reg [7:0] z2781_assgn2781;
    wire [7:0] z_x1_G256_newbasis1;
    wire [7:0] z_tempy2_G256_newbasis1;
    wire [7:0] z6443_assgn6443;
    reg [7:0] z6443_assgn64430;
    reg [7:0] z6443_assgn64431;
    reg [7:0] z6443_assgn64432;
    reg [7:0] z6443_assgn64433;
    reg [7:0] z6443_assgn64434;
    reg [7:0] z2785_assgn2785;
    wire [7:0] z_cond2_G256_newbasis1;
    wire [7:0] z_negCond2_G256_newbasis1;
    wire [7:0] z6449_assgn6449;
    reg [7:0] z6449_assgn64490;
    reg [7:0] z6449_assgn64491;
    reg [7:0] z6449_assgn64492;
    reg [7:0] z6449_assgn64493;
    reg [7:0] z6449_assgn64494;
    reg [7:0] z2789_assgn2789;
    wire [7:0] z_yxorb2_G256_newbasis1;
    wire [7:0] z_ny2_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond2_G256_newbasis1;
    wire [7:0] z_y2_G256_newbasis1;
    wire [7:0] z6459_assgn6459;
    reg [7:0] z6459_assgn64590;
    reg [7:0] z6459_assgn64591;
    reg [7:0] z6459_assgn64592;
    reg [7:0] z6459_assgn64593;
    reg [7:0] z6459_assgn64594;
    reg [7:0] z2797_assgn2797;
    wire [7:0] z_x2_G256_newbasis1;
    wire [7:0] z_tempy3_G256_newbasis1;
    wire [7:0] z6465_assgn6465;
    reg [7:0] z6465_assgn64650;
    reg [7:0] z6465_assgn64651;
    reg [7:0] z6465_assgn64652;
    reg [7:0] z6465_assgn64653;
    reg [7:0] z6465_assgn64654;
    reg [7:0] z2801_assgn2801;
    wire [7:0] z_cond3_G256_newbasis1;
    wire [7:0] z_negCond3_G256_newbasis1;
    wire [7:0] z6471_assgn6471;
    reg [7:0] z6471_assgn64710;
    reg [7:0] z6471_assgn64711;
    reg [7:0] z6471_assgn64712;
    reg [7:0] z6471_assgn64713;
    reg [7:0] z6471_assgn64714;
    reg [7:0] z2805_assgn2805;
    wire [7:0] z_yxorb3_G256_newbasis1;
    wire [7:0] z_ny3_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond3_G256_newbasis1;
    wire [7:0] z_y3_G256_newbasis1;
    wire [7:0] z6481_assgn6481;
    reg [7:0] z6481_assgn64810;
    reg [7:0] z6481_assgn64811;
    reg [7:0] z6481_assgn64812;
    reg [7:0] z6481_assgn64813;
    reg [7:0] z6481_assgn64814;
    reg [7:0] z2813_assgn2813;
    wire [7:0] z_x3_G256_newbasis1;
    wire [7:0] z_tempy4_G256_newbasis1;
    wire [7:0] z6487_assgn6487;
    reg [7:0] z6487_assgn64870;
    reg [7:0] z6487_assgn64871;
    reg [7:0] z6487_assgn64872;
    reg [7:0] z6487_assgn64873;
    reg [7:0] z6487_assgn64874;
    reg [7:0] z2817_assgn2817;
    wire [7:0] z_cond4_G256_newbasis1;
    wire [7:0] z_negCond4_G256_newbasis1;
    wire [7:0] z6493_assgn6493;
    reg [7:0] z6493_assgn64930;
    reg [7:0] z6493_assgn64931;
    reg [7:0] z6493_assgn64932;
    reg [7:0] z6493_assgn64933;
    reg [7:0] z6493_assgn64934;
    reg [7:0] z2821_assgn2821;
    wire [7:0] z_yxorb4_G256_newbasis1;
    wire [7:0] z_ny4_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond4_G256_newbasis1;
    wire [7:0] z_y4_G256_newbasis1;
    wire [7:0] z6503_assgn6503;
    reg [7:0] z6503_assgn65030;
    reg [7:0] z6503_assgn65031;
    reg [7:0] z6503_assgn65032;
    reg [7:0] z6503_assgn65033;
    reg [7:0] z6503_assgn65034;
    reg [7:0] z2829_assgn2829;
    wire [7:0] z_x4_G256_newbasis1;
    wire [7:0] z_tempy5_G256_newbasis1;
    wire [7:0] z6509_assgn6509;
    reg [7:0] z6509_assgn65090;
    reg [7:0] z6509_assgn65091;
    reg [7:0] z6509_assgn65092;
    reg [7:0] z6509_assgn65093;
    reg [7:0] z6509_assgn65094;
    reg [7:0] z2833_assgn2833;
    wire [7:0] z_cond5_G256_newbasis1;
    wire [7:0] z_negCond5_G256_newbasis1;
    wire [7:0] z6515_assgn6515;
    reg [7:0] z6515_assgn65150;
    reg [7:0] z6515_assgn65151;
    reg [7:0] z6515_assgn65152;
    reg [7:0] z6515_assgn65153;
    reg [7:0] z6515_assgn65154;
    reg [7:0] z2837_assgn2837;
    wire [7:0] z_yxorb5_G256_newbasis1;
    wire [7:0] z_ny5_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond5_G256_newbasis1;
    wire [7:0] z_y5_G256_newbasis1;
    wire [7:0] z6525_assgn6525;
    reg [7:0] z6525_assgn65250;
    reg [7:0] z6525_assgn65251;
    reg [7:0] z6525_assgn65252;
    reg [7:0] z6525_assgn65253;
    reg [7:0] z6525_assgn65254;
    reg [7:0] z2845_assgn2845;
    wire [7:0] z_x5_G256_newbasis1;
    wire [7:0] z_tempy6_G256_newbasis1;
    wire [7:0] z6531_assgn6531;
    reg [7:0] z6531_assgn65310;
    reg [7:0] z6531_assgn65311;
    reg [7:0] z6531_assgn65312;
    reg [7:0] z6531_assgn65313;
    reg [7:0] z6531_assgn65314;
    reg [7:0] z2849_assgn2849;
    wire [7:0] z_cond6_G256_newbasis1;
    wire [7:0] z_negCond6_G256_newbasis1;
    wire [7:0] z6537_assgn6537;
    reg [7:0] z6537_assgn65370;
    reg [7:0] z6537_assgn65371;
    reg [7:0] z6537_assgn65372;
    reg [7:0] z6537_assgn65373;
    reg [7:0] z6537_assgn65374;
    reg [7:0] z2853_assgn2853;
    wire [7:0] z_yxorb6_G256_newbasis1;
    wire [7:0] z_ny6_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond6_G256_newbasis1;
    wire [7:0] z_y6_G256_newbasis1;
    wire [7:0] z6547_assgn6547;
    reg [7:0] z6547_assgn65470;
    reg [7:0] z6547_assgn65471;
    reg [7:0] z6547_assgn65472;
    reg [7:0] z6547_assgn65473;
    reg [7:0] z6547_assgn65474;
    reg [7:0] z2861_assgn2861;
    wire [7:0] z_x6_G256_newbasis1;
    wire [7:0] z_tempy7_G256_newbasis1;
    wire [7:0] z6553_assgn6553;
    reg [7:0] z6553_assgn65530;
    reg [7:0] z6553_assgn65531;
    reg [7:0] z6553_assgn65532;
    reg [7:0] z6553_assgn65533;
    reg [7:0] z6553_assgn65534;
    reg [7:0] z2865_assgn2865;
    wire [7:0] z_cond7_G256_newbasis1;
    wire [7:0] z_negCond7_G256_newbasis1;
    wire [7:0] z6559_assgn6559;
    reg [7:0] z6559_assgn65590;
    reg [7:0] z6559_assgn65591;
    reg [7:0] z6559_assgn65592;
    reg [7:0] z6559_assgn65593;
    reg [7:0] z6559_assgn65594;
    reg [7:0] z2869_assgn2869;
    wire [7:0] z_yxorb7_G256_newbasis1;
    wire [7:0] z_ny7_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond7_G256_newbasis1;
    wire [7:0] z_y7_G256_newbasis1;
    wire [7:0] z6569_assgn6569;
    reg [7:0] z6569_assgn65690;
    reg [7:0] z6569_assgn65691;
    reg [7:0] z6569_assgn65692;
    reg [7:0] z6569_assgn65693;
    reg [7:0] z6569_assgn65694;
    reg [7:0] z2877_assgn2877;
    wire [7:0] z_x7_G256_newbasis1;
    wire [7:0] z_tempy8_G256_newbasis1;
    wire [7:0] z6575_assgn6575;
    reg [7:0] z6575_assgn65750;
    reg [7:0] z6575_assgn65751;
    reg [7:0] z6575_assgn65752;
    reg [7:0] z6575_assgn65753;
    reg [7:0] z6575_assgn65754;
    reg [7:0] z2881_assgn2881;
    wire [7:0] z_cond8_G256_newbasis1;
    wire [7:0] z_negCond8_G256_newbasis1;
    wire [7:0] z6581_assgn6581;
    reg [7:0] z6581_assgn65810;
    reg [7:0] z6581_assgn65811;
    reg [7:0] z6581_assgn65812;
    reg [7:0] z6581_assgn65813;
    reg [7:0] z6581_assgn65814;
    reg [7:0] z2885_assgn2885;
    wire [7:0] z_yxorb8_G256_newbasis1;
    wire [7:0] z_ny8_G256_newbasis1;
    wire [7:0] z_tempyIntoNegCond8_G256_newbasis1;
    wire [7:0] z_y8_G256_newbasis1;
    wire [7:0] z6591_assgn6591;
    reg [7:0] z6591_assgn65910;
    reg [7:0] z6591_assgn65911;
    reg [7:0] z6591_assgn65912;
    reg [7:0] z6591_assgn65913;
    reg [7:0] z6591_assgn65914;
    reg [7:0] z2893_assgn2893;
    wire [7:0] z_x8_G256_newbasis1;
    wire [7:0] t7;
    wire [7:0] z6597_assgn6597;
    reg [7:0] z6597_assgn65970;
    reg [7:0] z6597_assgn65971;
    reg [7:0] z6597_assgn65972;
    reg [7:0] z6597_assgn65973;
    reg [7:0] z6597_assgn65974;
    reg [7:0] z2897_assgn2897;

    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign r6_inp = r6;
    assign r7_inp = r7;
    assign r8_inp = r8;
    assign r9_inp = r9;
    assign r10_inp = r10;
    assign r11_inp = r11;
    assign r12_inp = r12;
    assign r13_inp = r13;
    assign r14_inp = r14;
    assign r15_inp = r15;
    assign r16_inp = r16;
    assign r17_inp = r17;
    assign r18_inp = r18;
    assign r19_inp = r19;
    assign r20_inp = r20;
    assign r21_inp = r21;
    assign r22_inp = r22;
    assign r23_inp = r23;
    assign r24_inp = r24;
    assign r25_inp = r25;
    assign r26_inp = r26;
    assign r27_inp = r27;
    assign r28_inp = r28;
    assign r29_inp = r29;
    assign r30_inp = r30;
    assign r31_inp = r31;
    assign r32_inp = r32;
    assign r33_inp = r33;
    assign r34_inp = r34;
    assign r35_inp = r35;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempyIntoNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempyIntoNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempyIntoNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempyIntoNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempyIntoNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempyIntoNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempyIntoNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempyIntoNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0);
    assign z3153_assgn3153 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempyIntoNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempyIntoNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempyIntoNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempyIntoNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempyIntoNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempyIntoNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempyIntoNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempyIntoNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempyIntoNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempyIntoNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempyIntoNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempyIntoNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempyIntoNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempyIntoNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempyIntoNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempyIntoNegCond8_G256_newbasis0);
    assign z3285_assgn3285 = (z_x7_G256_newbasis0 >> dec_1_inp);
    assign t3 = z_y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a1_0_G256_inv0 = (t3 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a1xorb1_G256_inv0 = (a1_G256_inv0 ^ b1_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul0_G256_inv0 = (r5_inp % dec_16_inp);
    assign r60_G16_mul0_G256_inv0 = (r6_inp % dec_16_inp);
    assign r70_G16_mul0_G256_inv0 = (r7_inp % dec_16_inp);
    assign r80_G16_mul0_G256_inv0 = (r8_inp % dec_16_inp);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ d1_G4_mul0_G16_mul0_G256_inv0);
    assign r0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 = !axorb_0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0 = !axorb_1_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign u1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign v0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign v1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign p0_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0_reg & cxord_0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0_reg & v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0_reg & cxord_1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc20_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0_reg & v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 = !a0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0 = !a1_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign u1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign v0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign v1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign p0_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0_reg & c0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0_reg & v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0_reg & c1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc21_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0_reg & v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul0_G256_inv0);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 = !b0_G4_mul0_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0 = !b1_G4_mul0_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign u1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign v0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (d0_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign v1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (d1_G4_mul0_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign p0_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0_reg & d0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0_reg & v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul0_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign p2_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0_reg & d1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_hpc22_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0_reg & v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul0_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul0_G256_inv0);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign z3583_assgn3583 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << z683_assgn683);
    assign z3587_assgn3587 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << z685_assgn685);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign z3595_assgn3595 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z691_assgn691);
    assign z3599_assgn3599 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z693_assgn693);
    assign z3603_assgn3603 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> z695_assgn695);
    assign z3607_assgn3607 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> z697_assgn697);
    assign z3611_assgn3611 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & z699_assgn699);
    assign z3615_assgn3615 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z701_assgn701);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign z3627_assgn3627 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << z711_assgn711);
    assign z3631_assgn3631 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << z713_assgn713);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ d1_G4_mul1_G16_mul0_G256_inv0);
    assign r0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 = !axorb_0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0 = !axorb_1_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign u1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign v0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (cxord_0_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign v1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (cxord_1_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign p0_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0_reg & cxord_0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0_reg & v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0_reg & cxord_1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc20_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0_reg & v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 = !a0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0 = !a1_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign u1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign v0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign v1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign p0_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0_reg & c0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0_reg & v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0_reg & c1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc21_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0_reg & v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 = !b0_G4_mul1_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0 = !b1_G4_mul1_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign u1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign v0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (d0_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign v1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (d1_G4_mul1_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign p0_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0_reg & d0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0_reg & v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul1_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign p2_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0_reg & d1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_hpc22_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0_reg & v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul1_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul0_G256_inv0);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign z3775_assgn3775 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << z855_assgn855);
    assign z3779_assgn3779 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << z857_assgn857);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r60_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r70_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r80_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ d1_G4_mul2_G16_mul0_G256_inv0);
    assign r0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 = !axorb_0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0 = !axorb_1_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign u1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign v0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (cxord_0_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign v1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (cxord_1_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign p0_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0_reg & cxord_0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0_reg & v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc20_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0_reg & cxord_1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc20_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0_reg & v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc20_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul0_G256_inv0);
    assign r0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 = !a0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0 = !a1_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign u1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign v0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign v1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign p0_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0_reg & c0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0_reg & v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc21_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0_reg & c1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc21_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0_reg & v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc21_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul0_G256_inv0);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign r0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 = !b0_G4_mul2_G16_mul0_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0 = !b1_G4_mul2_G16_mul0_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign u1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg & r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign v0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (d0_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign v1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (d1_G4_mul2_G16_mul0_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign p0_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0_reg & d0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0_reg & v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p01_hpc22_G4_mul2_G16_mul0_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign p2_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0_reg & d1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_hpc22_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0_reg & v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p23_hpc22_G4_mul2_G16_mul0_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign z3927_assgn3927 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << z1003_assgn1003);
    assign z3931_assgn3931 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << z1005_assgn1005);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign z3943_assgn3943 = dec_2_inp;
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << z1015_assgn1015);
    assign z3947_assgn3947 = dec_2_inp;
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << z1017_assgn1017);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign z3955_assgn3955 = c0_G256_inv0;
    assign c0xord0_G256_inv0 = (z1024_assgn1024 ^ d0_G256_inv0);
    assign z3959_assgn3959 = c1_G256_inv0;
    assign c1xord1_G256_inv0 = (z1026_assgn1026 ^ d1_G256_inv0);
    assign r00_G16_inv0_G256_inv0 = (r9_inp % dec_16_inp);
    assign r10_G16_inv0_G256_inv0 = (r10_inp % dec_16_inp);
    assign r20_G16_inv0_G256_inv0 = (r11_inp % dec_16_inp);
    assign r30_G16_inv0_G256_inv0 = (r12_inp % dec_16_inp);
    assign r40_G16_inv0_G256_inv0 = (r13_inp % dec_16_inp);
    assign r50_G16_inv0_G256_inv0 = (r14_inp % dec_16_inp);
    assign r60_G16_inv0_G256_inv0 = (r15_inp % dec_16_inp);
    assign r70_G16_inv0_G256_inv0 = (r16_inp % dec_16_inp);
    assign r80_G16_inv0_G256_inv0 = (r17_inp % dec_16_inp);
    assign z3981_assgn3981 = dec_12_inp;
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & z1045_assgn1045);
    assign z3985_assgn3985 = dec_12_inp;
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1047_assgn1047);
    assign z3989_assgn3989 = dec_2_inp;
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> z1049_assgn1049);
    assign z3993_assgn3993 = dec_2_inp;
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> z1051_assgn1051);
    assign z3997_assgn3997 = dec_3_inp;
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & z1053_assgn1053);
    assign z4001_assgn4001 = dec_3_inp;
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1055_assgn1055);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a1xorb1_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 ^ b1_G16_inv0_G256_inv0);
    assign z4009_assgn4009 = dec_2_inp;
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1061_assgn1061);
    assign z4013_assgn4013 = dec_2_inp;
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1063_assgn1063);
    assign z4017_assgn4017 = dec_1_inp;
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> z1065_assgn1065);
    assign z4021_assgn4021 = dec_1_inp;
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> z1067_assgn1067);
    assign z4025_assgn4025 = dec_1_inp;
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & z1069_assgn1069);
    assign z4029_assgn4029 = dec_1_inp;
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1071_assgn1071);
    assign z4033_assgn4033 = dec_1_inp;
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << z1073_assgn1073);
    assign z4037_assgn4037 = dec_1_inp;
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << z1075_assgn1075);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign z4045_assgn4045 = dec_2_inp;
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1081_assgn1081);
    assign z4049_assgn4049 = dec_2_inp;
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1083_assgn1083);
    assign z4053_assgn4053 = dec_1_inp;
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1085_assgn1085);
    assign z4057_assgn4057 = dec_1_inp;
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1087_assgn1087);
    assign z4061_assgn4061 = dec_1_inp;
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & z1089_assgn1089);
    assign z4065_assgn4065 = dec_1_inp;
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1091_assgn1091);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign z4077_assgn4077 = dec_1_inp;
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << z1101_assgn1101);
    assign z4081_assgn4081 = dec_1_inp;
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << z1103_assgn1103);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4095_assgn4095 = dec_2_inp;
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1115_assgn1115);
    assign z4099_assgn4099 = dec_2_inp;
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1117_assgn1117);
    assign z4103_assgn4103 = dec_1_inp;
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> z1119_assgn1119);
    assign z4107_assgn4107 = dec_1_inp;
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> z1121_assgn1121);
    assign z4111_assgn4111 = dec_1_inp;
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1123_assgn1123);
    assign z4115_assgn4115 = dec_1_inp;
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1125_assgn1125);
    assign z4119_assgn4119 = dec_2_inp;
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1127_assgn1127);
    assign z4123_assgn4123 = dec_2_inp;
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1129_assgn1129);
    assign z4127_assgn4127 = dec_1_inp;
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> z1131_assgn1131);
    assign z4131_assgn4131 = dec_1_inp;
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> z1133_assgn1133);
    assign z4135_assgn4135 = dec_1_inp;
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1135_assgn1135);
    assign z4139_assgn4139 = dec_1_inp;
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1137_assgn1137);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ d1_G4_mul3_G16_inv0_G256_inv0);
    assign r0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 = !axorb_0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 = !axorb_1_G4_mul3_G16_inv0_G256_inv0;
    assign z4157_assgn4157 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 & z1153_assgn1153);
    assign z4161_assgn4161 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul3_G16_inv0_G256_inv0 & z1155_assgn1155);
    assign z4165_assgn4165 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign v0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (cxord_0_G4_mul3_G16_inv0_G256_inv0 ^ z1157_assgn1157);
    assign z4169_assgn4169 = r0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign v1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (cxord_1_G4_mul3_G16_inv0_G256_inv0 ^ z1159_assgn1159);
    assign p0_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0_reg & cxord_0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0_reg & v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4177_assgn4177 = u0_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign p01_hpc20_G4_mul3_G16_inv0_G256_inv0 = (z1166_assgn1166 ^ p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul3_G16_inv0_G256_inv0);
    assign p2_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0_reg & cxord_1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_hpc20_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0_reg & v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4187_assgn4187 = u1_hpc20_G4_mul3_G16_inv0_G256_inv0;
    assign p23_hpc20_G4_mul3_G16_inv0_G256_inv0 = (z1174_assgn1174 ^ p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul3_G16_inv0_G256_inv0);
    assign r0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 = !a0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 = !a1_G4_mul3_G16_inv0_G256_inv0;
    assign z4199_assgn4199 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 & z1183_assgn1183);
    assign z4203_assgn4203 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul3_G16_inv0_G256_inv0 & z1185_assgn1185);
    assign z4207_assgn4207 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ z1187_assgn1187);
    assign z4211_assgn4211 = r0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ z1189_assgn1189);
    assign p0_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0_reg & c0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0_reg & v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4219_assgn4219 = u0_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign p01_hpc21_G4_mul3_G16_inv0_G256_inv0 = (z1196_assgn1196 ^ p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul3_G16_inv0_G256_inv0);
    assign p2_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0_reg & c1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_hpc21_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0_reg & v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4229_assgn4229 = u1_hpc21_G4_mul3_G16_inv0_G256_inv0;
    assign p23_hpc21_G4_mul3_G16_inv0_G256_inv0 = (z1204_assgn1204 ^ p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul3_G16_inv0_G256_inv0);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign r0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 = !b0_G4_mul3_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 = !b1_G4_mul3_G16_inv0_G256_inv0;
    assign z4245_assgn4245 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 & z1217_assgn1217);
    assign z4249_assgn4249 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul3_G16_inv0_G256_inv0 & z1219_assgn1219);
    assign z4253_assgn4253 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (d0_G4_mul3_G16_inv0_G256_inv0 ^ z1221_assgn1221);
    assign z4257_assgn4257 = r0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (d1_G4_mul3_G16_inv0_G256_inv0 ^ z1223_assgn1223);
    assign p0_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0_reg & d0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p1_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0_reg & v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4265_assgn4265 = u0_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign p01_hpc22_G4_mul3_G16_inv0_G256_inv0 = (z1230_assgn1230 ^ p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul3_G16_inv0_G256_inv0);
    assign p2_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0_reg & d1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p3_hpc22_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0_reg & v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z4275_assgn4275 = u1_hpc22_G4_mul3_G16_inv0_G256_inv0;
    assign p23_hpc22_G4_mul3_G16_inv0_G256_inv0 = (z1238_assgn1238 ^ p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul3_G16_inv0_G256_inv0);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign z4285_assgn4285 = dec_1_inp;
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << z1245_assgn1245);
    assign z4289_assgn4289 = dec_1_inp;
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << z1247_assgn1247);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign z4297_assgn4297 = c0_G16_inv0_G256_inv0;
    assign c0xord0_G16_inv0_G256_inv0 = (z1254_assgn1254 ^ d0_G16_inv0_G256_inv0);
    assign z4301_assgn4301 = c1_G16_inv0_G256_inv0;
    assign c1xord1_G16_inv0_G256_inv0 = (z1256_assgn1256 ^ d1_G16_inv0_G256_inv0);
    assign z4305_assgn4305 = dec_2_inp;
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1257_assgn1257);
    assign z4309_assgn4309 = dec_2_inp;
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1259_assgn1259);
    assign z4313_assgn4313 = dec_1_inp;
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> z1261_assgn1261);
    assign z4317_assgn4317 = dec_1_inp;
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> z1263_assgn1263);
    assign z4321_assgn4321 = dec_1_inp;
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & z1265_assgn1265);
    assign z4325_assgn4325 = dec_1_inp;
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1267_assgn1267);
    assign z4329_assgn4329 = dec_1_inp;
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << z1269_assgn1269);
    assign z4333_assgn4333 = dec_1_inp;
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << z1271_assgn1271);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4347_assgn4347 = dec_2_inp;
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1283_assgn1283);
    assign z4351_assgn4351 = dec_2_inp;
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1285_assgn1285);
    assign z4355_assgn4355 = dec_1_inp;
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> z1287_assgn1287);
    assign z4359_assgn4359 = dec_1_inp;
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> z1289_assgn1289);
    assign z4363_assgn4363 = dec_1_inp;
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1291_assgn1291);
    assign z4367_assgn4367 = dec_1_inp;
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1293_assgn1293);
    assign z4371_assgn4371 = dec_2_inp;
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1295_assgn1295);
    assign z4375_assgn4375 = dec_2_inp;
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1297_assgn1297);
    assign z4379_assgn4379 = dec_1_inp;
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> z1299_assgn1299);
    assign z4383_assgn4383 = dec_1_inp;
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> z1301_assgn1301);
    assign z4387_assgn4387 = dec_1_inp;
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & z1303_assgn1303);
    assign z4391_assgn4391 = dec_1_inp;
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1305_assgn1305);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ d1_G4_mul4_G16_inv0_G256_inv0);
    assign r0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 = !axorb_0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 = !axorb_1_G4_mul4_G16_inv0_G256_inv0;
    assign z4409_assgn4409 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 & z1321_assgn1321);
    assign z4413_assgn4413 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul4_G16_inv0_G256_inv0 & z1323_assgn1323);
    assign z4417_assgn4417 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign v0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (cxord_0_G4_mul4_G16_inv0_G256_inv0 ^ z1325_assgn1325);
    assign z4421_assgn4421 = r0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign v1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (cxord_1_G4_mul4_G16_inv0_G256_inv0 ^ z1327_assgn1327);
    assign z4425_assgn4425 = cxord_0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & z1329_assgn1329);
    assign z4429_assgn4429 = v1_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 & z1331_assgn1331);
    assign p01_hpc20_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul4_G16_inv0_G256_inv0);
    assign z4437_assgn4437 = cxord_1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & z1337_assgn1337);
    assign z4441_assgn4441 = v0_hpc20_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc20_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 & z1339_assgn1339);
    assign p23_hpc20_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul4_G16_inv0_G256_inv0);
    assign r0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 = !a0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 = !a1_G4_mul4_G16_inv0_G256_inv0;
    assign z4455_assgn4455 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 & z1351_assgn1351);
    assign z4459_assgn4459 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul4_G16_inv0_G256_inv0 & z1353_assgn1353);
    assign z4463_assgn4463 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ z1355_assgn1355);
    assign z4467_assgn4467 = r0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ z1357_assgn1357);
    assign z4471_assgn4471 = c0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & z1359_assgn1359);
    assign z4475_assgn4475 = v1_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 & z1361_assgn1361);
    assign p01_hpc21_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul4_G16_inv0_G256_inv0);
    assign z4483_assgn4483 = c1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & z1367_assgn1367);
    assign z4487_assgn4487 = v0_hpc21_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc21_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 & z1369_assgn1369);
    assign p23_hpc21_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul4_G16_inv0_G256_inv0);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign r0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 = !b0_G4_mul4_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 = !b1_G4_mul4_G16_inv0_G256_inv0;
    assign z4505_assgn4505 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 & z1385_assgn1385);
    assign z4509_assgn4509 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul4_G16_inv0_G256_inv0 & z1387_assgn1387);
    assign z4513_assgn4513 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (d0_G4_mul4_G16_inv0_G256_inv0 ^ z1389_assgn1389);
    assign z4517_assgn4517 = r0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (d1_G4_mul4_G16_inv0_G256_inv0 ^ z1391_assgn1391);
    assign z4521_assgn4521 = d0_G4_mul4_G16_inv0_G256_inv0;
    assign p0_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & z1393_assgn1393);
    assign z4525_assgn4525 = v1_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign p1_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 & z1395_assgn1395);
    assign p01_hpc22_G4_mul4_G16_inv0_G256_inv0 = (u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul4_G16_inv0_G256_inv0);
    assign z4533_assgn4533 = d1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & z1401_assgn1401);
    assign z4537_assgn4537 = v0_hpc22_G4_mul4_G16_inv0_G256_inv0;
    assign p3_hpc22_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 & z1403_assgn1403);
    assign p23_hpc22_G4_mul4_G16_inv0_G256_inv0 = (u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul4_G16_inv0_G256_inv0);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign z4549_assgn4549 = dec_1_inp;
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << z1413_assgn1413);
    assign z4553_assgn4553 = dec_1_inp;
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << z1415_assgn1415);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r60_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r70_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r80_G16_inv0_G256_inv0 % dec_4_inp);
    assign z4567_assgn4567 = dec_2_inp;
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1427_assgn1427);
    assign z4571_assgn4571 = dec_2_inp;
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1429_assgn1429);
    assign z4575_assgn4575 = dec_1_inp;
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> z1431_assgn1431);
    assign z4579_assgn4579 = dec_1_inp;
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> z1433_assgn1433);
    assign z4583_assgn4583 = dec_1_inp;
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & z1435_assgn1435);
    assign z4587_assgn4587 = dec_1_inp;
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1437_assgn1437);
    assign z4591_assgn4591 = dec_2_inp;
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1439_assgn1439);
    assign z4595_assgn4595 = dec_2_inp;
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1441_assgn1441);
    assign z4599_assgn4599 = dec_1_inp;
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> z1443_assgn1443);
    assign z4603_assgn4603 = dec_1_inp;
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> z1445_assgn1445);
    assign z4607_assgn4607 = dec_1_inp;
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & z1447_assgn1447);
    assign z4611_assgn4611 = dec_1_inp;
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1449_assgn1449);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ d1_G4_mul5_G16_inv0_G256_inv0);
    assign r0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 = !axorb_0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 = !axorb_1_G4_mul5_G16_inv0_G256_inv0;
    assign z4629_assgn4629 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 & z1465_assgn1465);
    assign z4633_assgn4633 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc20_G4_mul5_G16_inv0_G256_inv0 & z1467_assgn1467);
    assign z4637_assgn4637 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign v0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (cxord_0_G4_mul5_G16_inv0_G256_inv0 ^ z1469_assgn1469);
    assign z4641_assgn4641 = r0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign v1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (cxord_1_G4_mul5_G16_inv0_G256_inv0 ^ z1471_assgn1471);
    assign z4645_assgn4645 = cxord_0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & z1473_assgn1473);
    assign z4649_assgn4649 = v1_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 & z1475_assgn1475);
    assign p01_hpc20_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc20_G4_mul5_G16_inv0_G256_inv0);
    assign z4657_assgn4657 = cxord_1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & z1481_assgn1481);
    assign z4661_assgn4661 = v0_hpc20_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc20_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 & z1483_assgn1483);
    assign p23_hpc20_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc20_G4_mul5_G16_inv0_G256_inv0);
    assign r0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 = !a0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 = !a1_G4_mul5_G16_inv0_G256_inv0;
    assign z4675_assgn4675 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 & z1495_assgn1495);
    assign z4679_assgn4679 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc21_G4_mul5_G16_inv0_G256_inv0 & z1497_assgn1497);
    assign z4683_assgn4683 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign v0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ z1499_assgn1499);
    assign z4687_assgn4687 = r0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign v1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ z1501_assgn1501);
    assign z4691_assgn4691 = c0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & z1503_assgn1503);
    assign z4695_assgn4695 = v1_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 & z1505_assgn1505);
    assign p01_hpc21_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc21_G4_mul5_G16_inv0_G256_inv0);
    assign z4703_assgn4703 = c1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & z1511_assgn1511);
    assign z4707_assgn4707 = v0_hpc21_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc21_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 & z1513_assgn1513);
    assign p23_hpc21_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc21_G4_mul5_G16_inv0_G256_inv0);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign r0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 = !b0_G4_mul5_G16_inv0_G256_inv0;
    assign a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 = !b1_G4_mul5_G16_inv0_G256_inv0;
    assign z4725_assgn4725 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign u0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (a0_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 & z1529_assgn1529);
    assign z4729_assgn4729 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign u1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (a1_neg_hpc22_G4_mul5_G16_inv0_G256_inv0 & z1531_assgn1531);
    assign z4733_assgn4733 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign v0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (d0_G4_mul5_G16_inv0_G256_inv0 ^ z1533_assgn1533);
    assign z4737_assgn4737 = r0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign v1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (d1_G4_mul5_G16_inv0_G256_inv0 ^ z1535_assgn1535);
    assign z4741_assgn4741 = d0_G4_mul5_G16_inv0_G256_inv0;
    assign p0_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & z1537_assgn1537);
    assign z4745_assgn4745 = v1_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign p1_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 & z1539_assgn1539);
    assign p01_hpc22_G4_mul5_G16_inv0_G256_inv0 = (u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p01_hpc22_G4_mul5_G16_inv0_G256_inv0);
    assign z4753_assgn4753 = d1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & z1545_assgn1545);
    assign z4757_assgn4757 = v0_hpc22_G4_mul5_G16_inv0_G256_inv0;
    assign p3_hpc22_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 & z1547_assgn1547);
    assign p23_hpc22_G4_mul5_G16_inv0_G256_inv0 = (u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg ^ p23_hpc22_G4_mul5_G16_inv0_G256_inv0);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign z4769_assgn4769 = dec_1_inp;
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << z1557_assgn1557);
    assign z4773_assgn4773 = dec_1_inp;
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << z1559_assgn1559);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign z4781_assgn4781 = dec_2_inp;
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << z1565_assgn1565);
    assign z4785_assgn4785 = dec_2_inp;
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << z1567_assgn1567);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign r00_G16_mul1_G256_inv0 = (r18_inp % dec_16_inp);
    assign r10_G16_mul1_G256_inv0 = (r19_inp % dec_16_inp);
    assign r20_G16_mul1_G256_inv0 = (r20_inp % dec_16_inp);
    assign r30_G16_mul1_G256_inv0 = (r21_inp % dec_16_inp);
    assign r40_G16_mul1_G256_inv0 = (r22_inp % dec_16_inp);
    assign r50_G16_mul1_G256_inv0 = (r23_inp % dec_16_inp);
    assign r60_G16_mul1_G256_inv0 = (r24_inp % dec_16_inp);
    assign r70_G16_mul1_G256_inv0 = (r25_inp % dec_16_inp);
    assign r80_G16_mul1_G256_inv0 = (r26_inp % dec_16_inp);
    assign z4811_assgn4811 = dec_12_inp;
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1591_assgn1591);
    assign z4815_assgn4815 = dec_12_inp;
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1593_assgn1593);
    assign z4819_assgn4819 = dec_2_inp;
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> z1595_assgn1595);
    assign z4823_assgn4823 = dec_2_inp;
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> z1597_assgn1597);
    assign z4827_assgn4827 = dec_3_inp;
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & z1599_assgn1599);
    assign z4831_assgn4831 = dec_3_inp;
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1601_assgn1601);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign z4861_assgn4861 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1629_assgn1629);
    assign z4865_assgn4865 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1631_assgn1631);
    assign z4869_assgn4869 = dec_1_inp;
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> z1633_assgn1633);
    assign z4873_assgn4873 = dec_1_inp;
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> z1635_assgn1635);
    assign z4877_assgn4877 = dec_1_inp;
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & z1637_assgn1637);
    assign z4881_assgn4881 = dec_1_inp;
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1639_assgn1639);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ d1_G4_mul0_G16_mul1_G256_inv0);
    assign r0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 = !axorb_0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 = !axorb_1_G4_mul0_G16_mul1_G256_inv0;
    assign z4911_assgn4911 = r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 & z1667_assgn1667);
    assign z4915_assgn4915 = r0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul1_G256_inv0 & z1669_assgn1669);
    assign v0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign v1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign z4923_assgn4923 = cxord_0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1675_assgn1675);
    assign z4927_assgn4927 = v1_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 & z1677_assgn1677);
    assign p01_hpc20_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign z4935_assgn4935 = cxord_1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1683_assgn1683);
    assign z4939_assgn4939 = v0_hpc20_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc20_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 & z1685_assgn1685);
    assign p23_hpc20_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul1_G256_inv0);
    assign r0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 = !a0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 = !a1_G4_mul0_G16_mul1_G256_inv0;
    assign z4953_assgn4953 = r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 & z1697_assgn1697);
    assign z4957_assgn4957 = r0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul1_G256_inv0 & z1699_assgn1699);
    assign v0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign v1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign z4965_assgn4965 = c0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1705_assgn1705);
    assign z4969_assgn4969 = v1_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 & z1707_assgn1707);
    assign p01_hpc21_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign z4977_assgn4977 = c1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1713_assgn1713);
    assign z4981_assgn4981 = v0_hpc21_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc21_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 & z1715_assgn1715);
    assign p23_hpc21_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul1_G256_inv0);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign r0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 = !b0_G4_mul0_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 = !b1_G4_mul0_G16_mul1_G256_inv0;
    assign z4999_assgn4999 = r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 & z1731_assgn1731);
    assign z5003_assgn5003 = r0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul1_G256_inv0 & z1733_assgn1733);
    assign v0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (d0_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign v1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (d1_G4_mul0_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign z5011_assgn5011 = d0_G4_mul0_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1739_assgn1739);
    assign z5015_assgn5015 = v1_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign p1_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 & z1741_assgn1741);
    assign p01_hpc22_G4_mul0_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign z5023_assgn5023 = d1_G4_mul0_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1747_assgn1747);
    assign z5027_assgn5027 = v0_hpc22_G4_mul0_G16_mul1_G256_inv0;
    assign p3_hpc22_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 & z1749_assgn1749);
    assign p23_hpc22_G4_mul0_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul1_G256_inv0);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign z5039_assgn5039 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << z1759_assgn1759);
    assign z5043_assgn5043 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << z1761_assgn1761);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign z5051_assgn5051 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1767_assgn1767);
    assign z5055_assgn5055 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1769_assgn1769);
    assign z5059_assgn5059 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1771_assgn1771);
    assign z5063_assgn5063 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> z1773_assgn1773);
    assign z5067_assgn5067 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & z1775_assgn1775);
    assign z5071_assgn5071 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z1777_assgn1777);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z5083_assgn5083 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << z1787_assgn1787);
    assign z5087_assgn5087 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << z1789_assgn1789);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign z5101_assgn5101 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1801_assgn1801);
    assign z5105_assgn5105 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1803_assgn1803);
    assign z5109_assgn5109 = dec_1_inp;
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> z1805_assgn1805);
    assign z5113_assgn5113 = dec_1_inp;
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> z1807_assgn1807);
    assign z5117_assgn5117 = dec_1_inp;
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & z1809_assgn1809);
    assign z5121_assgn5121 = dec_1_inp;
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z1811_assgn1811);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ d1_G4_mul1_G16_mul1_G256_inv0);
    assign r0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 = !axorb_0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 = !axorb_1_G4_mul1_G16_mul1_G256_inv0;
    assign z5151_assgn5151 = r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 & z1839_assgn1839);
    assign z5155_assgn5155 = r0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul1_G256_inv0 & z1841_assgn1841);
    assign v0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (cxord_0_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign v1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (cxord_1_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign z5163_assgn5163 = cxord_0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1847_assgn1847);
    assign z5167_assgn5167 = v1_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 & z1849_assgn1849);
    assign p01_hpc20_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign z5175_assgn5175 = cxord_1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1855_assgn1855);
    assign z5179_assgn5179 = v0_hpc20_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc20_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 & z1857_assgn1857);
    assign p23_hpc20_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul1_G256_inv0);
    assign r0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 = !a0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 = !a1_G4_mul1_G16_mul1_G256_inv0;
    assign z5193_assgn5193 = r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 & z1869_assgn1869);
    assign z5197_assgn5197 = r0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul1_G256_inv0 & z1871_assgn1871);
    assign v0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign v1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign z5205_assgn5205 = c0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1877_assgn1877);
    assign z5209_assgn5209 = v1_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 & z1879_assgn1879);
    assign p01_hpc21_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign z5217_assgn5217 = c1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1885_assgn1885);
    assign z5221_assgn5221 = v0_hpc21_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc21_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 & z1887_assgn1887);
    assign p23_hpc21_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign r0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 = !b0_G4_mul1_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 = !b1_G4_mul1_G16_mul1_G256_inv0;
    assign z5239_assgn5239 = r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 & z1903_assgn1903);
    assign z5243_assgn5243 = r0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul1_G256_inv0 & z1905_assgn1905);
    assign v0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (d0_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign v1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (d1_G4_mul1_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign z5251_assgn5251 = d0_G4_mul1_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1911_assgn1911);
    assign z5255_assgn5255 = v1_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign p1_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 & z1913_assgn1913);
    assign p01_hpc22_G4_mul1_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign z5263_assgn5263 = d1_G4_mul1_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1919_assgn1919);
    assign z5267_assgn5267 = v0_hpc22_G4_mul1_G16_mul1_G256_inv0;
    assign p3_hpc22_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 & z1921_assgn1921);
    assign p23_hpc22_G4_mul1_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul1_G256_inv0);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign z5279_assgn5279 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << z1931_assgn1931);
    assign z5283_assgn5283 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << z1933_assgn1933);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r60_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r70_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r80_G16_mul1_G256_inv0 % dec_4_inp);
    assign z5301_assgn5301 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1949_assgn1949);
    assign z5305_assgn5305 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1951_assgn1951);
    assign z5309_assgn5309 = dec_1_inp;
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> z1953_assgn1953);
    assign z5313_assgn5313 = dec_1_inp;
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> z1955_assgn1955);
    assign z5317_assgn5317 = dec_1_inp;
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & z1957_assgn1957);
    assign z5321_assgn5321 = dec_1_inp;
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z1959_assgn1959);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ d1_G4_mul2_G16_mul1_G256_inv0);
    assign r0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 = !axorb_0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 = !axorb_1_G4_mul2_G16_mul1_G256_inv0;
    assign z5351_assgn5351 = r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 & z1987_assgn1987);
    assign z5355_assgn5355 = r0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul1_G256_inv0 & z1989_assgn1989);
    assign v0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (cxord_0_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign v1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (cxord_1_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign z5363_assgn5363 = cxord_0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z1995_assgn1995);
    assign z5367_assgn5367 = v1_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 & z1997_assgn1997);
    assign p01_hpc20_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign z5375_assgn5375 = cxord_1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z2003_assgn2003);
    assign z5379_assgn5379 = v0_hpc20_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc20_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 & z2005_assgn2005);
    assign p23_hpc20_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul1_G256_inv0);
    assign r0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 = !a0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 = !a1_G4_mul2_G16_mul1_G256_inv0;
    assign z5393_assgn5393 = r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 & z2017_assgn2017);
    assign z5397_assgn5397 = r0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul1_G256_inv0 & z2019_assgn2019);
    assign v0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign v1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign z5405_assgn5405 = c0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z2025_assgn2025);
    assign z5409_assgn5409 = v1_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 & z2027_assgn2027);
    assign p01_hpc21_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign z5417_assgn5417 = c1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z2033_assgn2033);
    assign z5421_assgn5421 = v0_hpc21_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc21_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 & z2035_assgn2035);
    assign p23_hpc21_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul1_G256_inv0);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign r0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 = !b0_G4_mul2_G16_mul1_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 = !b1_G4_mul2_G16_mul1_G256_inv0;
    assign z5439_assgn5439 = r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 & z2051_assgn2051);
    assign z5443_assgn5443 = r0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign u1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul1_G256_inv0 & z2053_assgn2053);
    assign v0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (d0_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign v1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (d1_G4_mul2_G16_mul1_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign z5451_assgn5451 = d0_G4_mul2_G16_mul1_G256_inv0;
    assign p0_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z2059_assgn2059);
    assign z5455_assgn5455 = v1_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign p1_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 & z2061_assgn2061);
    assign p01_hpc22_G4_mul2_G16_mul1_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign z5463_assgn5463 = d1_G4_mul2_G16_mul1_G256_inv0;
    assign p2_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z2067_assgn2067);
    assign z5467_assgn5467 = v0_hpc22_G4_mul2_G16_mul1_G256_inv0;
    assign p3_hpc22_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 & z2069_assgn2069);
    assign p23_hpc22_G4_mul2_G16_mul1_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign z5479_assgn5479 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << z2079_assgn2079);
    assign z5483_assgn5483 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << z2081_assgn2081);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign z5495_assgn5495 = dec_2_inp;
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << z2091_assgn2091);
    assign z5499_assgn5499 = dec_2_inp;
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << z2093_assgn2093);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign r00_G16_mul2_G256_inv0 = (r27_inp % dec_16_inp);
    assign r10_G16_mul2_G256_inv0 = (r28_inp % dec_16_inp);
    assign r20_G16_mul2_G256_inv0 = (r29_inp % dec_16_inp);
    assign r30_G16_mul2_G256_inv0 = (r30_inp % dec_16_inp);
    assign r40_G16_mul2_G256_inv0 = (r31_inp % dec_16_inp);
    assign r50_G16_mul2_G256_inv0 = (r32_inp % dec_16_inp);
    assign r60_G16_mul2_G256_inv0 = (r33_inp % dec_16_inp);
    assign r70_G16_mul2_G256_inv0 = (r34_inp % dec_16_inp);
    assign r80_G16_mul2_G256_inv0 = (r35_inp % dec_16_inp);
    assign z5525_assgn5525 = dec_12_inp;
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2117_assgn2117);
    assign z5529_assgn5529 = dec_12_inp;
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2119_assgn2119);
    assign z5533_assgn5533 = dec_2_inp;
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> z2121_assgn2121);
    assign z5537_assgn5537 = dec_2_inp;
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> z2123_assgn2123);
    assign z5541_assgn5541 = dec_3_inp;
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & z2125_assgn2125);
    assign z5545_assgn5545 = dec_3_inp;
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2127_assgn2127);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign z5575_assgn5575 = dec_2_inp;
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2155_assgn2155);
    assign z5579_assgn5579 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2157_assgn2157);
    assign z5583_assgn5583 = dec_1_inp;
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> z2159_assgn2159);
    assign z5587_assgn5587 = dec_1_inp;
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> z2161_assgn2161);
    assign z5591_assgn5591 = dec_1_inp;
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & z2163_assgn2163);
    assign z5595_assgn5595 = dec_1_inp;
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2165_assgn2165);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ d1_G4_mul0_G16_mul2_G256_inv0);
    assign r0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 = !axorb_0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 = !axorb_1_G4_mul0_G16_mul2_G256_inv0;
    assign z5625_assgn5625 = r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 & z2193_assgn2193);
    assign z5629_assgn5629 = r0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul0_G16_mul2_G256_inv0 & z2195_assgn2195);
    assign v0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign v1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign z5637_assgn5637 = cxord_0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z2201_assgn2201);
    assign z5641_assgn5641 = v1_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 & z2203_assgn2203);
    assign p01_hpc20_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign z5649_assgn5649 = cxord_1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z2209_assgn2209);
    assign z5653_assgn5653 = v0_hpc20_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc20_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 & z2211_assgn2211);
    assign p23_hpc20_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul0_G16_mul2_G256_inv0);
    assign r0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 = !a0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 = !a1_G4_mul0_G16_mul2_G256_inv0;
    assign z5667_assgn5667 = r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 & z2223_assgn2223);
    assign z5671_assgn5671 = r0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul0_G16_mul2_G256_inv0 & z2225_assgn2225);
    assign v0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign v1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign z5679_assgn5679 = c0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z2231_assgn2231);
    assign z5683_assgn5683 = v1_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 & z2233_assgn2233);
    assign p01_hpc21_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign z5691_assgn5691 = c1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z2239_assgn2239);
    assign z5695_assgn5695 = v0_hpc21_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc21_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 & z2241_assgn2241);
    assign p23_hpc21_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul0_G16_mul2_G256_inv0);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign r0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 = !b0_G4_mul0_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 = !b1_G4_mul0_G16_mul2_G256_inv0;
    assign z5713_assgn5713 = r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 & z2257_assgn2257);
    assign z5717_assgn5717 = r0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul0_G16_mul2_G256_inv0 & z2259_assgn2259);
    assign v0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (d0_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign v1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (d1_G4_mul0_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign z5725_assgn5725 = d0_G4_mul0_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z2265_assgn2265);
    assign z5729_assgn5729 = v1_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign p1_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 & z2267_assgn2267);
    assign p01_hpc22_G4_mul0_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign z5737_assgn5737 = d1_G4_mul0_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z2273_assgn2273);
    assign z5741_assgn5741 = v0_hpc22_G4_mul0_G16_mul2_G256_inv0;
    assign p3_hpc22_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 & z2275_assgn2275);
    assign p23_hpc22_G4_mul0_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul0_G16_mul2_G256_inv0);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign z5753_assgn5753 = dec_1_inp;
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << z2285_assgn2285);
    assign z5757_assgn5757 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << z2287_assgn2287);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign z5765_assgn5765 = dec_2_inp;
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2293_assgn2293);
    assign z5769_assgn5769 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2295_assgn2295);
    assign z5773_assgn5773 = dec_1_inp;
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2297_assgn2297);
    assign z5777_assgn5777 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2299_assgn2299);
    assign z5781_assgn5781 = dec_1_inp;
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & z2301_assgn2301);
    assign z5785_assgn5785 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2303_assgn2303);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z5797_assgn5797 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << z2313_assgn2313);
    assign z5801_assgn5801 = dec_1_inp;
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << z2315_assgn2315);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign z5815_assgn5815 = dec_2_inp;
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2327_assgn2327);
    assign z5819_assgn5819 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2329_assgn2329);
    assign z5823_assgn5823 = dec_1_inp;
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> z2331_assgn2331);
    assign z5827_assgn5827 = dec_1_inp;
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> z2333_assgn2333);
    assign z5831_assgn5831 = dec_1_inp;
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & z2335_assgn2335);
    assign z5835_assgn5835 = dec_1_inp;
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2337_assgn2337);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ d1_G4_mul1_G16_mul2_G256_inv0);
    assign r0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 = !axorb_0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 = !axorb_1_G4_mul1_G16_mul2_G256_inv0;
    assign z5865_assgn5865 = r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 & z2365_assgn2365);
    assign z5869_assgn5869 = r0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul1_G16_mul2_G256_inv0 & z2367_assgn2367);
    assign v0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (cxord_0_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign v1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (cxord_1_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign z5877_assgn5877 = cxord_0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2373_assgn2373);
    assign z5881_assgn5881 = v1_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 & z2375_assgn2375);
    assign p01_hpc20_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign z5889_assgn5889 = cxord_1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2381_assgn2381);
    assign z5893_assgn5893 = v0_hpc20_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc20_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 & z2383_assgn2383);
    assign p23_hpc20_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul1_G16_mul2_G256_inv0);
    assign r0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 = !a0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 = !a1_G4_mul1_G16_mul2_G256_inv0;
    assign z5907_assgn5907 = r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 & z2395_assgn2395);
    assign z5911_assgn5911 = r0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul1_G16_mul2_G256_inv0 & z2397_assgn2397);
    assign v0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign v1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign z5919_assgn5919 = c0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2403_assgn2403);
    assign z5923_assgn5923 = v1_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 & z2405_assgn2405);
    assign p01_hpc21_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign z5931_assgn5931 = c1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2411_assgn2411);
    assign z5935_assgn5935 = v0_hpc21_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc21_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 & z2413_assgn2413);
    assign p23_hpc21_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign r0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 = !b0_G4_mul1_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 = !b1_G4_mul1_G16_mul2_G256_inv0;
    assign z5953_assgn5953 = r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 & z2429_assgn2429);
    assign z5957_assgn5957 = r0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul1_G16_mul2_G256_inv0 & z2431_assgn2431);
    assign v0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (d0_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign v1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (d1_G4_mul1_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign z5965_assgn5965 = d0_G4_mul1_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2437_assgn2437);
    assign z5969_assgn5969 = v1_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign p1_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 & z2439_assgn2439);
    assign p01_hpc22_G4_mul1_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign z5977_assgn5977 = d1_G4_mul1_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2445_assgn2445);
    assign z5981_assgn5981 = v0_hpc22_G4_mul1_G16_mul2_G256_inv0;
    assign p3_hpc22_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 & z2447_assgn2447);
    assign p23_hpc22_G4_mul1_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul1_G16_mul2_G256_inv0);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign z5993_assgn5993 = dec_1_inp;
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << z2457_assgn2457);
    assign z5997_assgn5997 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << z2459_assgn2459);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r60_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r70_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r80_G16_mul2_G256_inv0 % dec_4_inp);
    assign z6015_assgn6015 = dec_2_inp;
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2475_assgn2475);
    assign z6019_assgn6019 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2477_assgn2477);
    assign z6023_assgn6023 = dec_1_inp;
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> z2479_assgn2479);
    assign z6027_assgn6027 = dec_1_inp;
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> z2481_assgn2481);
    assign z6031_assgn6031 = dec_1_inp;
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & z2483_assgn2483);
    assign z6035_assgn6035 = dec_1_inp;
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z2485_assgn2485);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ d1_G4_mul2_G16_mul2_G256_inv0);
    assign r0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 = !axorb_0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 = !axorb_1_G4_mul2_G16_mul2_G256_inv0;
    assign z6065_assgn6065 = r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 & z2513_assgn2513);
    assign z6069_assgn6069 = r0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc20_G4_mul2_G16_mul2_G256_inv0 & z2515_assgn2515);
    assign v0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (cxord_0_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign v1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (cxord_1_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign z6077_assgn6077 = cxord_0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2521_assgn2521);
    assign z6081_assgn6081 = v1_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 & z2523_assgn2523);
    assign p01_hpc20_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign z6089_assgn6089 = cxord_1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2529_assgn2529);
    assign z6093_assgn6093 = v0_hpc20_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc20_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 & z2531_assgn2531);
    assign p23_hpc20_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc20_G4_mul2_G16_mul2_G256_inv0);
    assign r0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 = !a0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 = !a1_G4_mul2_G16_mul2_G256_inv0;
    assign z6107_assgn6107 = r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 & z2543_assgn2543);
    assign z6111_assgn6111 = r0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc21_G4_mul2_G16_mul2_G256_inv0 & z2545_assgn2545);
    assign v0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign v1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign z6119_assgn6119 = c0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2551_assgn2551);
    assign z6123_assgn6123 = v1_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 & z2553_assgn2553);
    assign p01_hpc21_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign z6131_assgn6131 = c1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2559_assgn2559);
    assign z6135_assgn6135 = v0_hpc21_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc21_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 & z2561_assgn2561);
    assign p23_hpc21_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc21_G4_mul2_G16_mul2_G256_inv0);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign r0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 = !b0_G4_mul2_G16_mul2_G256_inv0;
    assign a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 = !b1_G4_mul2_G16_mul2_G256_inv0;
    assign z6153_assgn6153 = r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign u0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (a0_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 & z2577_assgn2577);
    assign z6157_assgn6157 = r0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign u1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (a1_neg_hpc22_G4_mul2_G16_mul2_G256_inv0 & z2579_assgn2579);
    assign v0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (d0_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign v1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (d1_G4_mul2_G16_mul2_G256_inv0 ^ r0_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign z6165_assgn6165 = d0_G4_mul2_G16_mul2_G256_inv0;
    assign p0_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2585_assgn2585);
    assign z6169_assgn6169 = v1_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign p1_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 & z2587_assgn2587);
    assign p01_hpc22_G4_mul2_G16_mul2_G256_inv0 = (u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p01_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign z6177_assgn6177 = d1_G4_mul2_G16_mul2_G256_inv0;
    assign p2_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2593_assgn2593);
    assign z6181_assgn6181 = v0_hpc22_G4_mul2_G16_mul2_G256_inv0;
    assign p3_hpc22_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 & z2595_assgn2595);
    assign p23_hpc22_G4_mul2_G16_mul2_G256_inv0 = (u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg ^ p23_hpc22_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign z6193_assgn6193 = dec_1_inp;
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << z2605_assgn2605);
    assign z6197_assgn6197 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << z2607_assgn2607);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign z6209_assgn6209 = dec_2_inp;
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << z2617_assgn2617);
    assign z6213_assgn6213 = dec_2_inp;
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << z2619_assgn2619);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign z6221_assgn6221 = dec_4_inp;
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << z2625_assgn2625);
    assign z6225_assgn6225 = dec_4_inp;
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << z2627_assgn2627);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign z6237_assgn6237 = dec_1_inp;
    assign cond1_G256_newbasis1 = (t4 & z2637_assgn2637);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign z6245_assgn6245 = yxorb1_G256_newbasis1;
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * z2643_assgn2643);
    assign z6249_assgn6249 = tempy1_G256_newbasis1;
    assign tempyIntoNegCond1_G256_newbasis1 = (z2646_assgn2646 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1);
    assign z6255_assgn6255 = dec_1_inp;
    assign x1_G256_newbasis1 = (t4 >> z2649_assgn2649);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign z6261_assgn6261 = dec_1_inp;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & z2653_assgn2653);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign z6267_assgn6267 = dec_3_inp;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ z2657_assgn2657);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempyIntoNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1);
    assign z6277_assgn6277 = dec_1_inp;
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> z2665_assgn2665);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign z6283_assgn6283 = dec_1_inp;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & z2669_assgn2669);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign z6289_assgn6289 = dec_4_inp;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ z2673_assgn2673);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempyIntoNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1);
    assign z6299_assgn6299 = dec_1_inp;
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> z2681_assgn2681);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign z6305_assgn6305 = dec_1_inp;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & z2685_assgn2685);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign z6311_assgn6311 = dec_220_inp;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ z2689_assgn2689);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempyIntoNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1);
    assign z6321_assgn6321 = dec_1_inp;
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> z2697_assgn2697);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign z6327_assgn6327 = dec_1_inp;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & z2701_assgn2701);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign z6333_assgn6333 = dec_11_inp;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ z2705_assgn2705);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempyIntoNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1);
    assign z6343_assgn6343 = dec_1_inp;
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> z2713_assgn2713);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign z6349_assgn6349 = dec_1_inp;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & z2717_assgn2717);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign z6355_assgn6355 = dec_158_inp;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ z2721_assgn2721);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempyIntoNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1);
    assign z6365_assgn6365 = dec_1_inp;
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> z2729_assgn2729);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign z6371_assgn6371 = dec_1_inp;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & z2733_assgn2733);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign z6377_assgn6377 = dec_45_inp;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ z2737_assgn2737);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempyIntoNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1);
    assign z6387_assgn6387 = dec_1_inp;
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> z2745_assgn2745);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign z6393_assgn6393 = dec_1_inp;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & z2749_assgn2749);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign z6399_assgn6399 = dec_88_inp;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ z2753_assgn2753);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempyIntoNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1);
    assign z6409_assgn6409 = dec_1_inp;
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> z2761_assgn2761);
    assign t6 = y8_G256_newbasis1;
    assign z_y_G256_newbasis1 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z6419_assgn6419 = dec_1_inp;
    assign z_cond1_G256_newbasis1 = (t5 & z2769_assgn2769);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z6427_assgn6427 = z_yxorb1_G256_newbasis1;
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z2775_assgn2775);
    assign z6431_assgn6431 = z_tempy1_G256_newbasis1;
    assign z_tempyIntoNegCond1_G256_newbasis1 = (z2778_assgn2778 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempyIntoNegCond1_G256_newbasis1);
    assign z6437_assgn6437 = dec_1_inp;
    assign z_x1_G256_newbasis1 = (t5 >> z2781_assgn2781);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z6443_assgn6443 = dec_1_inp;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & z2785_assgn2785);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z6449_assgn6449 = dec_3_inp;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ z2789_assgn2789);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempyIntoNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempyIntoNegCond2_G256_newbasis1);
    assign z6459_assgn6459 = dec_1_inp;
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> z2797_assgn2797);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z6465_assgn6465 = dec_1_inp;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & z2801_assgn2801);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z6471_assgn6471 = dec_4_inp;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ z2805_assgn2805);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempyIntoNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempyIntoNegCond3_G256_newbasis1);
    assign z6481_assgn6481 = dec_1_inp;
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> z2813_assgn2813);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z6487_assgn6487 = dec_1_inp;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & z2817_assgn2817);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z6493_assgn6493 = dec_220_inp;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ z2821_assgn2821);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempyIntoNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempyIntoNegCond4_G256_newbasis1);
    assign z6503_assgn6503 = dec_1_inp;
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> z2829_assgn2829);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z6509_assgn6509 = dec_1_inp;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & z2833_assgn2833);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z6515_assgn6515 = dec_11_inp;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ z2837_assgn2837);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempyIntoNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempyIntoNegCond5_G256_newbasis1);
    assign z6525_assgn6525 = dec_1_inp;
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> z2845_assgn2845);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z6531_assgn6531 = dec_1_inp;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & z2849_assgn2849);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z6537_assgn6537 = dec_158_inp;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ z2853_assgn2853);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempyIntoNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempyIntoNegCond6_G256_newbasis1);
    assign z6547_assgn6547 = dec_1_inp;
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> z2861_assgn2861);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z6553_assgn6553 = dec_1_inp;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & z2865_assgn2865);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z6559_assgn6559 = dec_45_inp;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ z2869_assgn2869);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempyIntoNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempyIntoNegCond7_G256_newbasis1);
    assign z6569_assgn6569 = dec_1_inp;
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> z2877_assgn2877);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z6575_assgn6575 = dec_1_inp;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & z2881_assgn2881);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z6581_assgn6581 = dec_88_inp;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ z2885_assgn2885);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempyIntoNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempyIntoNegCond8_G256_newbasis1);
    assign z6591_assgn6591 = dec_1_inp;
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> z2893_assgn2893);
    assign t7 = z_y8_G256_newbasis1;
    assign z6597_assgn6597 = dec_99_inp;

    always @(posedge clk) begin
        z3153_assgn31530 <= z3153_assgn3153;
        z3153_assgn31531 <= z3153_assgn31530;
        z3153_assgn31532 <= z3153_assgn31531;
        z3153_assgn31533 <= z3153_assgn31532;
        z3153_assgn31534 <= z3153_assgn31533;
        x8_G256_newbasis0 <= z3153_assgn31534;
        z3285_assgn32850 <= z3285_assgn3285;
        z3285_assgn32851 <= z3285_assgn32850;
        z3285_assgn32852 <= z3285_assgn32851;
        z3285_assgn32853 <= z3285_assgn32852;
        z3285_assgn32854 <= z3285_assgn32853;
        z_x8_G256_newbasis0 <= z3285_assgn32854;
        a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= a0_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= a1_neg_hpc20_G4_mul0_G16_mul0_G256_inv0;
        axorb_0_G4_mul0_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul0_G16_mul0_G256_inv0;
        cxord_0_G4_mul0_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul0_G16_mul0_G256_inv0;
        v1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        axorb_1_G4_mul0_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul0_G16_mul0_G256_inv0;
        cxord_1_G4_mul0_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul0_G16_mul0_G256_inv0;
        v0_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul0_G256_inv0;
        a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= a0_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
        r0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= a1_neg_hpc21_G4_mul0_G16_mul0_G256_inv0;
        a0_G4_mul0_G16_mul0_G256_inv0_reg <= a0_G4_mul0_G16_mul0_G256_inv0;
        c0_G4_mul0_G16_mul0_G256_inv0_reg <= c0_G4_mul0_G16_mul0_G256_inv0;
        v1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        a1_G4_mul0_G16_mul0_G256_inv0_reg <= a1_G4_mul0_G16_mul0_G256_inv0;
        c1_G4_mul0_G16_mul0_G256_inv0_reg <= c1_G4_mul0_G16_mul0_G256_inv0;
        v0_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul0_G256_inv0;
        a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= a0_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
        r0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= a1_neg_hpc22_G4_mul0_G16_mul0_G256_inv0;
        b0_G4_mul0_G16_mul0_G256_inv0_reg <= b0_G4_mul0_G16_mul0_G256_inv0;
        d0_G4_mul0_G16_mul0_G256_inv0_reg <= d0_G4_mul0_G16_mul0_G256_inv0;
        v1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        b1_G4_mul0_G16_mul0_G256_inv0_reg <= b1_G4_mul0_G16_mul0_G256_inv0;
        d1_G4_mul0_G16_mul0_G256_inv0_reg <= d1_G4_mul0_G16_mul0_G256_inv0;
        v0_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul0_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul0_G256_inv0;
        z3583_assgn35830 <= z3583_assgn3583;
        z683_assgn683 <= z3583_assgn35830;
        z3587_assgn35870 <= z3587_assgn3587;
        z685_assgn685 <= z3587_assgn35870;
        z3595_assgn35950 <= z3595_assgn3595;
        z691_assgn691 <= z3595_assgn35950;
        z3599_assgn35990 <= z3599_assgn3599;
        z693_assgn693 <= z3599_assgn35990;
        z3603_assgn36030 <= z3603_assgn3603;
        z695_assgn695 <= z3603_assgn36030;
        z3607_assgn36070 <= z3607_assgn3607;
        z697_assgn697 <= z3607_assgn36070;
        z3611_assgn36110 <= z3611_assgn3611;
        z699_assgn699 <= z3611_assgn36110;
        z3615_assgn36150 <= z3615_assgn3615;
        z701_assgn701 <= z3615_assgn36150;
        z3627_assgn36270 <= z3627_assgn3627;
        z711_assgn711 <= z3627_assgn36270;
        z3631_assgn36310 <= z3631_assgn3631;
        z713_assgn713 <= z3631_assgn36310;
        a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= a0_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= a1_neg_hpc20_G4_mul1_G16_mul0_G256_inv0;
        axorb_0_G4_mul1_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul1_G16_mul0_G256_inv0;
        cxord_0_G4_mul1_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul1_G16_mul0_G256_inv0;
        v1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        axorb_1_G4_mul1_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul1_G16_mul0_G256_inv0;
        cxord_1_G4_mul1_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul1_G16_mul0_G256_inv0;
        v0_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul0_G256_inv0;
        a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= a0_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
        r0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= a1_neg_hpc21_G4_mul1_G16_mul0_G256_inv0;
        a0_G4_mul1_G16_mul0_G256_inv0_reg <= a0_G4_mul1_G16_mul0_G256_inv0;
        c0_G4_mul1_G16_mul0_G256_inv0_reg <= c0_G4_mul1_G16_mul0_G256_inv0;
        v1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        a1_G4_mul1_G16_mul0_G256_inv0_reg <= a1_G4_mul1_G16_mul0_G256_inv0;
        c1_G4_mul1_G16_mul0_G256_inv0_reg <= c1_G4_mul1_G16_mul0_G256_inv0;
        v0_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul0_G256_inv0;
        a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= a0_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
        r0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= a1_neg_hpc22_G4_mul1_G16_mul0_G256_inv0;
        b0_G4_mul1_G16_mul0_G256_inv0_reg <= b0_G4_mul1_G16_mul0_G256_inv0;
        d0_G4_mul1_G16_mul0_G256_inv0_reg <= d0_G4_mul1_G16_mul0_G256_inv0;
        v1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        b1_G4_mul1_G16_mul0_G256_inv0_reg <= b1_G4_mul1_G16_mul0_G256_inv0;
        d1_G4_mul1_G16_mul0_G256_inv0_reg <= d1_G4_mul1_G16_mul0_G256_inv0;
        v0_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul1_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul0_G256_inv0;
        z3775_assgn37750 <= z3775_assgn3775;
        z855_assgn855 <= z3775_assgn37750;
        z3779_assgn37790 <= z3779_assgn3779;
        z857_assgn857 <= z3779_assgn37790;
        a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= a0_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
        r0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= a1_neg_hpc20_G4_mul2_G16_mul0_G256_inv0;
        axorb_0_G4_mul2_G16_mul0_G256_inv0_reg <= axorb_0_G4_mul2_G16_mul0_G256_inv0;
        cxord_0_G4_mul2_G16_mul0_G256_inv0_reg <= cxord_0_G4_mul2_G16_mul0_G256_inv0;
        v1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        axorb_1_G4_mul2_G16_mul0_G256_inv0_reg <= axorb_1_G4_mul2_G16_mul0_G256_inv0;
        cxord_1_G4_mul2_G16_mul0_G256_inv0_reg <= cxord_1_G4_mul2_G16_mul0_G256_inv0;
        v0_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc20_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul0_G256_inv0;
        a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= a0_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
        r0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= a1_neg_hpc21_G4_mul2_G16_mul0_G256_inv0;
        a0_G4_mul2_G16_mul0_G256_inv0_reg <= a0_G4_mul2_G16_mul0_G256_inv0;
        c0_G4_mul2_G16_mul0_G256_inv0_reg <= c0_G4_mul2_G16_mul0_G256_inv0;
        v1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        a1_G4_mul2_G16_mul0_G256_inv0_reg <= a1_G4_mul2_G16_mul0_G256_inv0;
        c1_G4_mul2_G16_mul0_G256_inv0_reg <= c1_G4_mul2_G16_mul0_G256_inv0;
        v0_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc21_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul0_G256_inv0;
        a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= a0_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
        r0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= r0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= a1_neg_hpc22_G4_mul2_G16_mul0_G256_inv0;
        b0_G4_mul2_G16_mul0_G256_inv0_reg <= b0_G4_mul2_G16_mul0_G256_inv0;
        d0_G4_mul2_G16_mul0_G256_inv0_reg <= d0_G4_mul2_G16_mul0_G256_inv0;
        v1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= v1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        u0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        b1_G4_mul2_G16_mul0_G256_inv0_reg <= b1_G4_mul2_G16_mul0_G256_inv0;
        d1_G4_mul2_G16_mul0_G256_inv0_reg <= d1_G4_mul2_G16_mul0_G256_inv0;
        v0_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= v0_hpc22_G4_mul2_G16_mul0_G256_inv0;
        u1_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul0_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul0_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul0_G256_inv0;
        z3927_assgn39270 <= z3927_assgn3927;
        z1003_assgn1003 <= z3927_assgn39270;
        z3931_assgn39310 <= z3931_assgn3931;
        z1005_assgn1005 <= z3931_assgn39310;
        z3943_assgn39430 <= z3943_assgn3943;
        z1015_assgn1015 <= z3943_assgn39430;
        z3947_assgn39470 <= z3947_assgn3947;
        z1017_assgn1017 <= z3947_assgn39470;
        z3955_assgn39550 <= z3955_assgn3955;
        z1024_assgn1024 <= z3955_assgn39550;
        z3959_assgn39590 <= z3959_assgn3959;
        z1026_assgn1026 <= z3959_assgn39590;
        z3981_assgn39810 <= z3981_assgn3981;
        z1045_assgn1045 <= z3981_assgn39810;
        z3985_assgn39850 <= z3985_assgn3985;
        z1047_assgn1047 <= z3985_assgn39850;
        z3989_assgn39890 <= z3989_assgn3989;
        z1049_assgn1049 <= z3989_assgn39890;
        z3993_assgn39930 <= z3993_assgn3993;
        z1051_assgn1051 <= z3993_assgn39930;
        z3997_assgn39970 <= z3997_assgn3997;
        z1053_assgn1053 <= z3997_assgn39970;
        z4001_assgn40010 <= z4001_assgn4001;
        z1055_assgn1055 <= z4001_assgn40010;
        z4009_assgn40090 <= z4009_assgn4009;
        z1061_assgn1061 <= z4009_assgn40090;
        z4013_assgn40130 <= z4013_assgn4013;
        z1063_assgn1063 <= z4013_assgn40130;
        z4017_assgn40170 <= z4017_assgn4017;
        z1065_assgn1065 <= z4017_assgn40170;
        z4021_assgn40210 <= z4021_assgn4021;
        z1067_assgn1067 <= z4021_assgn40210;
        z4025_assgn40250 <= z4025_assgn4025;
        z1069_assgn1069 <= z4025_assgn40250;
        z4029_assgn40290 <= z4029_assgn4029;
        z1071_assgn1071 <= z4029_assgn40290;
        z4033_assgn40330 <= z4033_assgn4033;
        z1073_assgn1073 <= z4033_assgn40330;
        z4037_assgn40370 <= z4037_assgn4037;
        z1075_assgn1075 <= z4037_assgn40370;
        z4045_assgn40450 <= z4045_assgn4045;
        z1081_assgn1081 <= z4045_assgn40450;
        z4049_assgn40490 <= z4049_assgn4049;
        z1083_assgn1083 <= z4049_assgn40490;
        z4053_assgn40530 <= z4053_assgn4053;
        z1085_assgn1085 <= z4053_assgn40530;
        z4057_assgn40570 <= z4057_assgn4057;
        z1087_assgn1087 <= z4057_assgn40570;
        z4061_assgn40610 <= z4061_assgn4061;
        z1089_assgn1089 <= z4061_assgn40610;
        z4065_assgn40650 <= z4065_assgn4065;
        z1091_assgn1091 <= z4065_assgn40650;
        z4077_assgn40770 <= z4077_assgn4077;
        z1101_assgn1101 <= z4077_assgn40770;
        z4081_assgn40810 <= z4081_assgn4081;
        z1103_assgn1103 <= z4081_assgn40810;
        z4095_assgn40950 <= z4095_assgn4095;
        z1115_assgn1115 <= z4095_assgn40950;
        z4099_assgn40990 <= z4099_assgn4099;
        z1117_assgn1117 <= z4099_assgn40990;
        z4103_assgn41030 <= z4103_assgn4103;
        z1119_assgn1119 <= z4103_assgn41030;
        z4107_assgn41070 <= z4107_assgn4107;
        z1121_assgn1121 <= z4107_assgn41070;
        z4111_assgn41110 <= z4111_assgn4111;
        z1123_assgn1123 <= z4111_assgn41110;
        z4115_assgn41150 <= z4115_assgn4115;
        z1125_assgn1125 <= z4115_assgn41150;
        z4119_assgn41190 <= z4119_assgn4119;
        z1127_assgn1127 <= z4119_assgn41190;
        z4123_assgn41230 <= z4123_assgn4123;
        z1129_assgn1129 <= z4123_assgn41230;
        z4127_assgn41270 <= z4127_assgn4127;
        z1131_assgn1131 <= z4127_assgn41270;
        z4131_assgn41310 <= z4131_assgn4131;
        z1133_assgn1133 <= z4131_assgn41310;
        z4135_assgn41350 <= z4135_assgn4135;
        z1135_assgn1135 <= z4135_assgn41350;
        z4139_assgn41390 <= z4139_assgn4139;
        z1137_assgn1137 <= z4139_assgn41390;
        z4157_assgn41570 <= z4157_assgn4157;
        z1153_assgn1153 <= z4157_assgn41570;
        z4161_assgn41610 <= z4161_assgn4161;
        z1155_assgn1155 <= z4161_assgn41610;
        z4165_assgn41650 <= z4165_assgn4165;
        z1157_assgn1157 <= z4165_assgn41650;
        z4169_assgn41690 <= z4169_assgn4169;
        z1159_assgn1159 <= z4169_assgn41690;
        axorb_0_G4_mul3_G16_inv0_G256_inv0_reg <= axorb_0_G4_mul3_G16_inv0_G256_inv0;
        cxord_0_G4_mul3_G16_inv0_G256_inv0_reg <= cxord_0_G4_mul3_G16_inv0_G256_inv0;
        v1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc20_G4_mul3_G16_inv0_G256_inv0;
        z4177_assgn41770 <= z4177_assgn4177;
        z1166_assgn1166 <= z4177_assgn41770;
        p1_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        axorb_1_G4_mul3_G16_inv0_G256_inv0_reg <= axorb_1_G4_mul3_G16_inv0_G256_inv0;
        cxord_1_G4_mul3_G16_inv0_G256_inv0_reg <= cxord_1_G4_mul3_G16_inv0_G256_inv0;
        v0_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc20_G4_mul3_G16_inv0_G256_inv0;
        z4187_assgn41870 <= z4187_assgn4187;
        z1174_assgn1174 <= z4187_assgn41870;
        p3_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul3_G16_inv0_G256_inv0;
        z4199_assgn41990 <= z4199_assgn4199;
        z1183_assgn1183 <= z4199_assgn41990;
        z4203_assgn42030 <= z4203_assgn4203;
        z1185_assgn1185 <= z4203_assgn42030;
        z4207_assgn42070 <= z4207_assgn4207;
        z1187_assgn1187 <= z4207_assgn42070;
        z4211_assgn42110 <= z4211_assgn4211;
        z1189_assgn1189 <= z4211_assgn42110;
        a0_G4_mul3_G16_inv0_G256_inv0_reg <= a0_G4_mul3_G16_inv0_G256_inv0;
        c0_G4_mul3_G16_inv0_G256_inv0_reg <= c0_G4_mul3_G16_inv0_G256_inv0;
        v1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4219_assgn42190 <= z4219_assgn4219;
        z1196_assgn1196 <= z4219_assgn42190;
        p1_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        a1_G4_mul3_G16_inv0_G256_inv0_reg <= a1_G4_mul3_G16_inv0_G256_inv0;
        c1_G4_mul3_G16_inv0_G256_inv0_reg <= c1_G4_mul3_G16_inv0_G256_inv0;
        v0_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4229_assgn42290 <= z4229_assgn4229;
        z1204_assgn1204 <= z4229_assgn42290;
        p3_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul3_G16_inv0_G256_inv0;
        z4245_assgn42450 <= z4245_assgn4245;
        z1217_assgn1217 <= z4245_assgn42450;
        z4249_assgn42490 <= z4249_assgn4249;
        z1219_assgn1219 <= z4249_assgn42490;
        z4253_assgn42530 <= z4253_assgn4253;
        z1221_assgn1221 <= z4253_assgn42530;
        z4257_assgn42570 <= z4257_assgn4257;
        z1223_assgn1223 <= z4257_assgn42570;
        b0_G4_mul3_G16_inv0_G256_inv0_reg <= b0_G4_mul3_G16_inv0_G256_inv0;
        d0_G4_mul3_G16_inv0_G256_inv0_reg <= d0_G4_mul3_G16_inv0_G256_inv0;
        v1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= v1_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4265_assgn42650 <= z4265_assgn4265;
        z1230_assgn1230 <= z4265_assgn42650;
        p1_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        b1_G4_mul3_G16_inv0_G256_inv0_reg <= b1_G4_mul3_G16_inv0_G256_inv0;
        d1_G4_mul3_G16_inv0_G256_inv0_reg <= d1_G4_mul3_G16_inv0_G256_inv0;
        v0_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= v0_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4275_assgn42750 <= z4275_assgn4275;
        z1238_assgn1238 <= z4275_assgn42750;
        p3_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul3_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul3_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul3_G16_inv0_G256_inv0;
        z4285_assgn42850 <= z4285_assgn4285;
        z4285_assgn42851 <= z4285_assgn42850;
        z4285_assgn42852 <= z4285_assgn42851;
        z1245_assgn1245 <= z4285_assgn42852;
        z4289_assgn42890 <= z4289_assgn4289;
        z4289_assgn42891 <= z4289_assgn42890;
        z4289_assgn42892 <= z4289_assgn42891;
        z1247_assgn1247 <= z4289_assgn42892;
        z4297_assgn42970 <= z4297_assgn4297;
        z1254_assgn1254 <= z4297_assgn42970;
        z4301_assgn43010 <= z4301_assgn4301;
        z1256_assgn1256 <= z4301_assgn43010;
        z4305_assgn43050 <= z4305_assgn4305;
        z4305_assgn43051 <= z4305_assgn43050;
        z4305_assgn43052 <= z4305_assgn43051;
        z1257_assgn1257 <= z4305_assgn43052;
        z4309_assgn43090 <= z4309_assgn4309;
        z4309_assgn43091 <= z4309_assgn43090;
        z4309_assgn43092 <= z4309_assgn43091;
        z1259_assgn1259 <= z4309_assgn43092;
        z4313_assgn43130 <= z4313_assgn4313;
        z4313_assgn43131 <= z4313_assgn43130;
        z4313_assgn43132 <= z4313_assgn43131;
        z1261_assgn1261 <= z4313_assgn43132;
        z4317_assgn43170 <= z4317_assgn4317;
        z4317_assgn43171 <= z4317_assgn43170;
        z4317_assgn43172 <= z4317_assgn43171;
        z1263_assgn1263 <= z4317_assgn43172;
        z4321_assgn43210 <= z4321_assgn4321;
        z4321_assgn43211 <= z4321_assgn43210;
        z4321_assgn43212 <= z4321_assgn43211;
        z1265_assgn1265 <= z4321_assgn43212;
        z4325_assgn43250 <= z4325_assgn4325;
        z4325_assgn43251 <= z4325_assgn43250;
        z4325_assgn43252 <= z4325_assgn43251;
        z1267_assgn1267 <= z4325_assgn43252;
        z4329_assgn43290 <= z4329_assgn4329;
        z4329_assgn43291 <= z4329_assgn43290;
        z4329_assgn43292 <= z4329_assgn43291;
        z1269_assgn1269 <= z4329_assgn43292;
        z4333_assgn43330 <= z4333_assgn4333;
        z4333_assgn43331 <= z4333_assgn43330;
        z4333_assgn43332 <= z4333_assgn43331;
        z1271_assgn1271 <= z4333_assgn43332;
        z4347_assgn43470 <= z4347_assgn4347;
        z4347_assgn43471 <= z4347_assgn43470;
        z4347_assgn43472 <= z4347_assgn43471;
        z1283_assgn1283 <= z4347_assgn43472;
        z4351_assgn43510 <= z4351_assgn4351;
        z4351_assgn43511 <= z4351_assgn43510;
        z4351_assgn43512 <= z4351_assgn43511;
        z1285_assgn1285 <= z4351_assgn43512;
        z4355_assgn43550 <= z4355_assgn4355;
        z4355_assgn43551 <= z4355_assgn43550;
        z4355_assgn43552 <= z4355_assgn43551;
        z1287_assgn1287 <= z4355_assgn43552;
        z4359_assgn43590 <= z4359_assgn4359;
        z4359_assgn43591 <= z4359_assgn43590;
        z4359_assgn43592 <= z4359_assgn43591;
        z1289_assgn1289 <= z4359_assgn43592;
        z4363_assgn43630 <= z4363_assgn4363;
        z4363_assgn43631 <= z4363_assgn43630;
        z4363_assgn43632 <= z4363_assgn43631;
        z1291_assgn1291 <= z4363_assgn43632;
        z4367_assgn43670 <= z4367_assgn4367;
        z4367_assgn43671 <= z4367_assgn43670;
        z4367_assgn43672 <= z4367_assgn43671;
        z1293_assgn1293 <= z4367_assgn43672;
        z4371_assgn43710 <= z4371_assgn4371;
        z1295_assgn1295 <= z4371_assgn43710;
        z4375_assgn43750 <= z4375_assgn4375;
        z1297_assgn1297 <= z4375_assgn43750;
        z4379_assgn43790 <= z4379_assgn4379;
        z1299_assgn1299 <= z4379_assgn43790;
        z4383_assgn43830 <= z4383_assgn4383;
        z1301_assgn1301 <= z4383_assgn43830;
        z4387_assgn43870 <= z4387_assgn4387;
        z1303_assgn1303 <= z4387_assgn43870;
        z4391_assgn43910 <= z4391_assgn4391;
        z1305_assgn1305 <= z4391_assgn43910;
        z4409_assgn44090 <= z4409_assgn4409;
        z4409_assgn44091 <= z4409_assgn44090;
        z4409_assgn44092 <= z4409_assgn44091;
        z1321_assgn1321 <= z4409_assgn44092;
        z4413_assgn44130 <= z4413_assgn4413;
        z4413_assgn44131 <= z4413_assgn44130;
        z4413_assgn44132 <= z4413_assgn44131;
        z1323_assgn1323 <= z4413_assgn44132;
        z4417_assgn44170 <= z4417_assgn4417;
        z1325_assgn1325 <= z4417_assgn44170;
        z4421_assgn44210 <= z4421_assgn4421;
        z1327_assgn1327 <= z4421_assgn44210;
        z4425_assgn44250 <= z4425_assgn4425;
        z1329_assgn1329 <= z4425_assgn44250;
        z4429_assgn44290 <= z4429_assgn4429;
        z1331_assgn1331 <= z4429_assgn44290;
        u0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul4_G16_inv0_G256_inv0;
        z4437_assgn44370 <= z4437_assgn4437;
        z1337_assgn1337 <= z4437_assgn44370;
        z4441_assgn44410 <= z4441_assgn4441;
        z1339_assgn1339 <= z4441_assgn44410;
        u1_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul4_G16_inv0_G256_inv0;
        z4455_assgn44550 <= z4455_assgn4455;
        z4455_assgn44551 <= z4455_assgn44550;
        z4455_assgn44552 <= z4455_assgn44551;
        z1351_assgn1351 <= z4455_assgn44552;
        z4459_assgn44590 <= z4459_assgn4459;
        z4459_assgn44591 <= z4459_assgn44590;
        z4459_assgn44592 <= z4459_assgn44591;
        z1353_assgn1353 <= z4459_assgn44592;
        z4463_assgn44630 <= z4463_assgn4463;
        z1355_assgn1355 <= z4463_assgn44630;
        z4467_assgn44670 <= z4467_assgn4467;
        z1357_assgn1357 <= z4467_assgn44670;
        z4471_assgn44710 <= z4471_assgn4471;
        z1359_assgn1359 <= z4471_assgn44710;
        z4475_assgn44750 <= z4475_assgn4475;
        z1361_assgn1361 <= z4475_assgn44750;
        u0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul4_G16_inv0_G256_inv0;
        z4483_assgn44830 <= z4483_assgn4483;
        z1367_assgn1367 <= z4483_assgn44830;
        z4487_assgn44870 <= z4487_assgn4487;
        z1369_assgn1369 <= z4487_assgn44870;
        u1_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul4_G16_inv0_G256_inv0;
        z4505_assgn45050 <= z4505_assgn4505;
        z4505_assgn45051 <= z4505_assgn45050;
        z4505_assgn45052 <= z4505_assgn45051;
        z1385_assgn1385 <= z4505_assgn45052;
        z4509_assgn45090 <= z4509_assgn4509;
        z4509_assgn45091 <= z4509_assgn45090;
        z4509_assgn45092 <= z4509_assgn45091;
        z1387_assgn1387 <= z4509_assgn45092;
        z4513_assgn45130 <= z4513_assgn4513;
        z1389_assgn1389 <= z4513_assgn45130;
        z4517_assgn45170 <= z4517_assgn4517;
        z1391_assgn1391 <= z4517_assgn45170;
        z4521_assgn45210 <= z4521_assgn4521;
        z1393_assgn1393 <= z4521_assgn45210;
        z4525_assgn45250 <= z4525_assgn4525;
        z1395_assgn1395 <= z4525_assgn45250;
        u0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= u0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul4_G16_inv0_G256_inv0;
        z4533_assgn45330 <= z4533_assgn4533;
        z1401_assgn1401 <= z4533_assgn45330;
        z4537_assgn45370 <= z4537_assgn4537;
        z1403_assgn1403 <= z4537_assgn45370;
        u1_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= u1_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p3_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul4_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul4_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul4_G16_inv0_G256_inv0;
        z4549_assgn45490 <= z4549_assgn4549;
        z4549_assgn45491 <= z4549_assgn45490;
        z4549_assgn45492 <= z4549_assgn45491;
        z4549_assgn45493 <= z4549_assgn45492;
        z1413_assgn1413 <= z4549_assgn45493;
        z4553_assgn45530 <= z4553_assgn4553;
        z4553_assgn45531 <= z4553_assgn45530;
        z4553_assgn45532 <= z4553_assgn45531;
        z4553_assgn45533 <= z4553_assgn45532;
        z1415_assgn1415 <= z4553_assgn45533;
        z4567_assgn45670 <= z4567_assgn4567;
        z4567_assgn45671 <= z4567_assgn45670;
        z4567_assgn45672 <= z4567_assgn45671;
        z1427_assgn1427 <= z4567_assgn45672;
        z4571_assgn45710 <= z4571_assgn4571;
        z4571_assgn45711 <= z4571_assgn45710;
        z4571_assgn45712 <= z4571_assgn45711;
        z1429_assgn1429 <= z4571_assgn45712;
        z4575_assgn45750 <= z4575_assgn4575;
        z4575_assgn45751 <= z4575_assgn45750;
        z4575_assgn45752 <= z4575_assgn45751;
        z1431_assgn1431 <= z4575_assgn45752;
        z4579_assgn45790 <= z4579_assgn4579;
        z4579_assgn45791 <= z4579_assgn45790;
        z4579_assgn45792 <= z4579_assgn45791;
        z1433_assgn1433 <= z4579_assgn45792;
        z4583_assgn45830 <= z4583_assgn4583;
        z4583_assgn45831 <= z4583_assgn45830;
        z4583_assgn45832 <= z4583_assgn45831;
        z1435_assgn1435 <= z4583_assgn45832;
        z4587_assgn45870 <= z4587_assgn4587;
        z4587_assgn45871 <= z4587_assgn45870;
        z4587_assgn45872 <= z4587_assgn45871;
        z1437_assgn1437 <= z4587_assgn45872;
        z4591_assgn45910 <= z4591_assgn4591;
        z1439_assgn1439 <= z4591_assgn45910;
        z4595_assgn45950 <= z4595_assgn4595;
        z1441_assgn1441 <= z4595_assgn45950;
        z4599_assgn45990 <= z4599_assgn4599;
        z1443_assgn1443 <= z4599_assgn45990;
        z4603_assgn46030 <= z4603_assgn4603;
        z1445_assgn1445 <= z4603_assgn46030;
        z4607_assgn46070 <= z4607_assgn4607;
        z1447_assgn1447 <= z4607_assgn46070;
        z4611_assgn46110 <= z4611_assgn4611;
        z1449_assgn1449 <= z4611_assgn46110;
        z4629_assgn46290 <= z4629_assgn4629;
        z4629_assgn46291 <= z4629_assgn46290;
        z4629_assgn46292 <= z4629_assgn46291;
        z1465_assgn1465 <= z4629_assgn46292;
        z4633_assgn46330 <= z4633_assgn4633;
        z4633_assgn46331 <= z4633_assgn46330;
        z4633_assgn46332 <= z4633_assgn46331;
        z1467_assgn1467 <= z4633_assgn46332;
        z4637_assgn46370 <= z4637_assgn4637;
        z1469_assgn1469 <= z4637_assgn46370;
        z4641_assgn46410 <= z4641_assgn4641;
        z1471_assgn1471 <= z4641_assgn46410;
        z4645_assgn46450 <= z4645_assgn4645;
        z1473_assgn1473 <= z4645_assgn46450;
        z4649_assgn46490 <= z4649_assgn4649;
        z1475_assgn1475 <= z4649_assgn46490;
        u0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc20_G4_mul5_G16_inv0_G256_inv0;
        z4657_assgn46570 <= z4657_assgn4657;
        z1481_assgn1481 <= z4657_assgn46570;
        z4661_assgn46610 <= z4661_assgn4661;
        z1483_assgn1483 <= z4661_assgn46610;
        u1_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc20_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc20_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc20_G4_mul5_G16_inv0_G256_inv0;
        z4675_assgn46750 <= z4675_assgn4675;
        z4675_assgn46751 <= z4675_assgn46750;
        z4675_assgn46752 <= z4675_assgn46751;
        z1495_assgn1495 <= z4675_assgn46752;
        z4679_assgn46790 <= z4679_assgn4679;
        z4679_assgn46791 <= z4679_assgn46790;
        z4679_assgn46792 <= z4679_assgn46791;
        z1497_assgn1497 <= z4679_assgn46792;
        z4683_assgn46830 <= z4683_assgn4683;
        z1499_assgn1499 <= z4683_assgn46830;
        z4687_assgn46870 <= z4687_assgn4687;
        z1501_assgn1501 <= z4687_assgn46870;
        z4691_assgn46910 <= z4691_assgn4691;
        z1503_assgn1503 <= z4691_assgn46910;
        z4695_assgn46950 <= z4695_assgn4695;
        z1505_assgn1505 <= z4695_assgn46950;
        u0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc21_G4_mul5_G16_inv0_G256_inv0;
        z4703_assgn47030 <= z4703_assgn4703;
        z1511_assgn1511 <= z4703_assgn47030;
        z4707_assgn47070 <= z4707_assgn4707;
        z1513_assgn1513 <= z4707_assgn47070;
        u1_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc21_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc21_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc21_G4_mul5_G16_inv0_G256_inv0;
        z4725_assgn47250 <= z4725_assgn4725;
        z4725_assgn47251 <= z4725_assgn47250;
        z4725_assgn47252 <= z4725_assgn47251;
        z1529_assgn1529 <= z4725_assgn47252;
        z4729_assgn47290 <= z4729_assgn4729;
        z4729_assgn47291 <= z4729_assgn47290;
        z4729_assgn47292 <= z4729_assgn47291;
        z1531_assgn1531 <= z4729_assgn47292;
        z4733_assgn47330 <= z4733_assgn4733;
        z1533_assgn1533 <= z4733_assgn47330;
        z4737_assgn47370 <= z4737_assgn4737;
        z1535_assgn1535 <= z4737_assgn47370;
        z4741_assgn47410 <= z4741_assgn4741;
        z1537_assgn1537 <= z4741_assgn47410;
        z4745_assgn47450 <= z4745_assgn4745;
        z1539_assgn1539 <= z4745_assgn47450;
        u0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= u0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p1_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p0_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p0_hpc22_G4_mul5_G16_inv0_G256_inv0;
        z4753_assgn47530 <= z4753_assgn4753;
        z1545_assgn1545 <= z4753_assgn47530;
        z4757_assgn47570 <= z4757_assgn4757;
        z1547_assgn1547 <= z4757_assgn47570;
        u1_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= u1_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p3_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p3_hpc22_G4_mul5_G16_inv0_G256_inv0;
        p2_hpc22_G4_mul5_G16_inv0_G256_inv0_reg <= p2_hpc22_G4_mul5_G16_inv0_G256_inv0;
        z4769_assgn47690 <= z4769_assgn4769;
        z4769_assgn47691 <= z4769_assgn47690;
        z4769_assgn47692 <= z4769_assgn47691;
        z4769_assgn47693 <= z4769_assgn47692;
        z1557_assgn1557 <= z4769_assgn47693;
        z4773_assgn47730 <= z4773_assgn4773;
        z4773_assgn47731 <= z4773_assgn47730;
        z4773_assgn47732 <= z4773_assgn47731;
        z4773_assgn47733 <= z4773_assgn47732;
        z1559_assgn1559 <= z4773_assgn47733;
        z4781_assgn47810 <= z4781_assgn4781;
        z4781_assgn47811 <= z4781_assgn47810;
        z4781_assgn47812 <= z4781_assgn47811;
        z4781_assgn47813 <= z4781_assgn47812;
        z1565_assgn1565 <= z4781_assgn47813;
        z4785_assgn47850 <= z4785_assgn4785;
        z4785_assgn47851 <= z4785_assgn47850;
        z4785_assgn47852 <= z4785_assgn47851;
        z4785_assgn47853 <= z4785_assgn47852;
        z1567_assgn1567 <= z4785_assgn47853;
        z4811_assgn48110 <= z4811_assgn4811;
        z4811_assgn48111 <= z4811_assgn48110;
        z4811_assgn48112 <= z4811_assgn48111;
        z4811_assgn48113 <= z4811_assgn48112;
        z1591_assgn1591 <= z4811_assgn48113;
        z4815_assgn48150 <= z4815_assgn4815;
        z4815_assgn48151 <= z4815_assgn48150;
        z4815_assgn48152 <= z4815_assgn48151;
        z4815_assgn48153 <= z4815_assgn48152;
        z1593_assgn1593 <= z4815_assgn48153;
        z4819_assgn48190 <= z4819_assgn4819;
        z4819_assgn48191 <= z4819_assgn48190;
        z4819_assgn48192 <= z4819_assgn48191;
        z4819_assgn48193 <= z4819_assgn48192;
        z1595_assgn1595 <= z4819_assgn48193;
        z4823_assgn48230 <= z4823_assgn4823;
        z4823_assgn48231 <= z4823_assgn48230;
        z4823_assgn48232 <= z4823_assgn48231;
        z4823_assgn48233 <= z4823_assgn48232;
        z1597_assgn1597 <= z4823_assgn48233;
        z4827_assgn48270 <= z4827_assgn4827;
        z4827_assgn48271 <= z4827_assgn48270;
        z4827_assgn48272 <= z4827_assgn48271;
        z4827_assgn48273 <= z4827_assgn48272;
        z1599_assgn1599 <= z4827_assgn48273;
        z4831_assgn48310 <= z4831_assgn4831;
        z4831_assgn48311 <= z4831_assgn48310;
        z4831_assgn48312 <= z4831_assgn48311;
        z4831_assgn48313 <= z4831_assgn48312;
        z1601_assgn1601 <= z4831_assgn48313;
        z4861_assgn48610 <= z4861_assgn4861;
        z4861_assgn48611 <= z4861_assgn48610;
        z4861_assgn48612 <= z4861_assgn48611;
        z4861_assgn48613 <= z4861_assgn48612;
        z1629_assgn1629 <= z4861_assgn48613;
        z4865_assgn48650 <= z4865_assgn4865;
        z4865_assgn48651 <= z4865_assgn48650;
        z4865_assgn48652 <= z4865_assgn48651;
        z4865_assgn48653 <= z4865_assgn48652;
        z1631_assgn1631 <= z4865_assgn48653;
        z4869_assgn48690 <= z4869_assgn4869;
        z4869_assgn48691 <= z4869_assgn48690;
        z4869_assgn48692 <= z4869_assgn48691;
        z4869_assgn48693 <= z4869_assgn48692;
        z1633_assgn1633 <= z4869_assgn48693;
        z4873_assgn48730 <= z4873_assgn4873;
        z4873_assgn48731 <= z4873_assgn48730;
        z4873_assgn48732 <= z4873_assgn48731;
        z4873_assgn48733 <= z4873_assgn48732;
        z1635_assgn1635 <= z4873_assgn48733;
        z4877_assgn48770 <= z4877_assgn4877;
        z4877_assgn48771 <= z4877_assgn48770;
        z4877_assgn48772 <= z4877_assgn48771;
        z4877_assgn48773 <= z4877_assgn48772;
        z1637_assgn1637 <= z4877_assgn48773;
        z4881_assgn48810 <= z4881_assgn4881;
        z4881_assgn48811 <= z4881_assgn48810;
        z4881_assgn48812 <= z4881_assgn48811;
        z4881_assgn48813 <= z4881_assgn48812;
        z1639_assgn1639 <= z4881_assgn48813;
        z4911_assgn49110 <= z4911_assgn4911;
        z4911_assgn49111 <= z4911_assgn49110;
        z4911_assgn49112 <= z4911_assgn49111;
        z4911_assgn49113 <= z4911_assgn49112;
        z1667_assgn1667 <= z4911_assgn49113;
        z4915_assgn49150 <= z4915_assgn4915;
        z4915_assgn49151 <= z4915_assgn49150;
        z4915_assgn49152 <= z4915_assgn49151;
        z4915_assgn49153 <= z4915_assgn49152;
        z1669_assgn1669 <= z4915_assgn49153;
        z4923_assgn49230 <= z4923_assgn4923;
        z4923_assgn49231 <= z4923_assgn49230;
        z4923_assgn49232 <= z4923_assgn49231;
        z4923_assgn49233 <= z4923_assgn49232;
        z1675_assgn1675 <= z4923_assgn49233;
        z4927_assgn49270 <= z4927_assgn4927;
        z4927_assgn49271 <= z4927_assgn49270;
        z4927_assgn49272 <= z4927_assgn49271;
        z4927_assgn49273 <= z4927_assgn49272;
        z1677_assgn1677 <= z4927_assgn49273;
        u0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul1_G256_inv0;
        z4935_assgn49350 <= z4935_assgn4935;
        z4935_assgn49351 <= z4935_assgn49350;
        z4935_assgn49352 <= z4935_assgn49351;
        z4935_assgn49353 <= z4935_assgn49352;
        z1683_assgn1683 <= z4935_assgn49353;
        z4939_assgn49390 <= z4939_assgn4939;
        z4939_assgn49391 <= z4939_assgn49390;
        z4939_assgn49392 <= z4939_assgn49391;
        z4939_assgn49393 <= z4939_assgn49392;
        z1685_assgn1685 <= z4939_assgn49393;
        u1_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul1_G256_inv0;
        z4953_assgn49530 <= z4953_assgn4953;
        z4953_assgn49531 <= z4953_assgn49530;
        z4953_assgn49532 <= z4953_assgn49531;
        z4953_assgn49533 <= z4953_assgn49532;
        z1697_assgn1697 <= z4953_assgn49533;
        z4957_assgn49570 <= z4957_assgn4957;
        z4957_assgn49571 <= z4957_assgn49570;
        z4957_assgn49572 <= z4957_assgn49571;
        z4957_assgn49573 <= z4957_assgn49572;
        z1699_assgn1699 <= z4957_assgn49573;
        z4965_assgn49650 <= z4965_assgn4965;
        z4965_assgn49651 <= z4965_assgn49650;
        z4965_assgn49652 <= z4965_assgn49651;
        z4965_assgn49653 <= z4965_assgn49652;
        z1705_assgn1705 <= z4965_assgn49653;
        z4969_assgn49690 <= z4969_assgn4969;
        z4969_assgn49691 <= z4969_assgn49690;
        z4969_assgn49692 <= z4969_assgn49691;
        z4969_assgn49693 <= z4969_assgn49692;
        z1707_assgn1707 <= z4969_assgn49693;
        u0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul1_G256_inv0;
        z4977_assgn49770 <= z4977_assgn4977;
        z4977_assgn49771 <= z4977_assgn49770;
        z4977_assgn49772 <= z4977_assgn49771;
        z4977_assgn49773 <= z4977_assgn49772;
        z1713_assgn1713 <= z4977_assgn49773;
        z4981_assgn49810 <= z4981_assgn4981;
        z4981_assgn49811 <= z4981_assgn49810;
        z4981_assgn49812 <= z4981_assgn49811;
        z4981_assgn49813 <= z4981_assgn49812;
        z1715_assgn1715 <= z4981_assgn49813;
        u1_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul1_G256_inv0;
        z4999_assgn49990 <= z4999_assgn4999;
        z4999_assgn49991 <= z4999_assgn49990;
        z4999_assgn49992 <= z4999_assgn49991;
        z4999_assgn49993 <= z4999_assgn49992;
        z1731_assgn1731 <= z4999_assgn49993;
        z5003_assgn50030 <= z5003_assgn5003;
        z5003_assgn50031 <= z5003_assgn50030;
        z5003_assgn50032 <= z5003_assgn50031;
        z5003_assgn50033 <= z5003_assgn50032;
        z1733_assgn1733 <= z5003_assgn50033;
        z5011_assgn50110 <= z5011_assgn5011;
        z5011_assgn50111 <= z5011_assgn50110;
        z5011_assgn50112 <= z5011_assgn50111;
        z5011_assgn50113 <= z5011_assgn50112;
        z1739_assgn1739 <= z5011_assgn50113;
        z5015_assgn50150 <= z5015_assgn5015;
        z5015_assgn50151 <= z5015_assgn50150;
        z5015_assgn50152 <= z5015_assgn50151;
        z5015_assgn50153 <= z5015_assgn50152;
        z1741_assgn1741 <= z5015_assgn50153;
        u0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul1_G256_inv0;
        z5023_assgn50230 <= z5023_assgn5023;
        z5023_assgn50231 <= z5023_assgn50230;
        z5023_assgn50232 <= z5023_assgn50231;
        z5023_assgn50233 <= z5023_assgn50232;
        z1747_assgn1747 <= z5023_assgn50233;
        z5027_assgn50270 <= z5027_assgn5027;
        z5027_assgn50271 <= z5027_assgn50270;
        z5027_assgn50272 <= z5027_assgn50271;
        z5027_assgn50273 <= z5027_assgn50272;
        z1749_assgn1749 <= z5027_assgn50273;
        u1_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul1_G256_inv0;
        z5039_assgn50390 <= z5039_assgn5039;
        z5039_assgn50391 <= z5039_assgn50390;
        z5039_assgn50392 <= z5039_assgn50391;
        z5039_assgn50393 <= z5039_assgn50392;
        z5039_assgn50394 <= z5039_assgn50393;
        z1759_assgn1759 <= z5039_assgn50394;
        z5043_assgn50430 <= z5043_assgn5043;
        z5043_assgn50431 <= z5043_assgn50430;
        z5043_assgn50432 <= z5043_assgn50431;
        z5043_assgn50433 <= z5043_assgn50432;
        z5043_assgn50434 <= z5043_assgn50433;
        z1761_assgn1761 <= z5043_assgn50434;
        z5051_assgn50510 <= z5051_assgn5051;
        z5051_assgn50511 <= z5051_assgn50510;
        z5051_assgn50512 <= z5051_assgn50511;
        z5051_assgn50513 <= z5051_assgn50512;
        z5051_assgn50514 <= z5051_assgn50513;
        z1767_assgn1767 <= z5051_assgn50514;
        z5055_assgn50550 <= z5055_assgn5055;
        z5055_assgn50551 <= z5055_assgn50550;
        z5055_assgn50552 <= z5055_assgn50551;
        z5055_assgn50553 <= z5055_assgn50552;
        z5055_assgn50554 <= z5055_assgn50553;
        z1769_assgn1769 <= z5055_assgn50554;
        z5059_assgn50590 <= z5059_assgn5059;
        z5059_assgn50591 <= z5059_assgn50590;
        z5059_assgn50592 <= z5059_assgn50591;
        z5059_assgn50593 <= z5059_assgn50592;
        z5059_assgn50594 <= z5059_assgn50593;
        z1771_assgn1771 <= z5059_assgn50594;
        z5063_assgn50630 <= z5063_assgn5063;
        z5063_assgn50631 <= z5063_assgn50630;
        z5063_assgn50632 <= z5063_assgn50631;
        z5063_assgn50633 <= z5063_assgn50632;
        z5063_assgn50634 <= z5063_assgn50633;
        z1773_assgn1773 <= z5063_assgn50634;
        z5067_assgn50670 <= z5067_assgn5067;
        z5067_assgn50671 <= z5067_assgn50670;
        z5067_assgn50672 <= z5067_assgn50671;
        z5067_assgn50673 <= z5067_assgn50672;
        z5067_assgn50674 <= z5067_assgn50673;
        z1775_assgn1775 <= z5067_assgn50674;
        z5071_assgn50710 <= z5071_assgn5071;
        z5071_assgn50711 <= z5071_assgn50710;
        z5071_assgn50712 <= z5071_assgn50711;
        z5071_assgn50713 <= z5071_assgn50712;
        z5071_assgn50714 <= z5071_assgn50713;
        z1777_assgn1777 <= z5071_assgn50714;
        z5083_assgn50830 <= z5083_assgn5083;
        z5083_assgn50831 <= z5083_assgn50830;
        z5083_assgn50832 <= z5083_assgn50831;
        z5083_assgn50833 <= z5083_assgn50832;
        z5083_assgn50834 <= z5083_assgn50833;
        z1787_assgn1787 <= z5083_assgn50834;
        z5087_assgn50870 <= z5087_assgn5087;
        z5087_assgn50871 <= z5087_assgn50870;
        z5087_assgn50872 <= z5087_assgn50871;
        z5087_assgn50873 <= z5087_assgn50872;
        z5087_assgn50874 <= z5087_assgn50873;
        z1789_assgn1789 <= z5087_assgn50874;
        z5101_assgn51010 <= z5101_assgn5101;
        z5101_assgn51011 <= z5101_assgn51010;
        z5101_assgn51012 <= z5101_assgn51011;
        z5101_assgn51013 <= z5101_assgn51012;
        z1801_assgn1801 <= z5101_assgn51013;
        z5105_assgn51050 <= z5105_assgn5105;
        z5105_assgn51051 <= z5105_assgn51050;
        z5105_assgn51052 <= z5105_assgn51051;
        z5105_assgn51053 <= z5105_assgn51052;
        z1803_assgn1803 <= z5105_assgn51053;
        z5109_assgn51090 <= z5109_assgn5109;
        z5109_assgn51091 <= z5109_assgn51090;
        z5109_assgn51092 <= z5109_assgn51091;
        z5109_assgn51093 <= z5109_assgn51092;
        z1805_assgn1805 <= z5109_assgn51093;
        z5113_assgn51130 <= z5113_assgn5113;
        z5113_assgn51131 <= z5113_assgn51130;
        z5113_assgn51132 <= z5113_assgn51131;
        z5113_assgn51133 <= z5113_assgn51132;
        z1807_assgn1807 <= z5113_assgn51133;
        z5117_assgn51170 <= z5117_assgn5117;
        z5117_assgn51171 <= z5117_assgn51170;
        z5117_assgn51172 <= z5117_assgn51171;
        z5117_assgn51173 <= z5117_assgn51172;
        z1809_assgn1809 <= z5117_assgn51173;
        z5121_assgn51210 <= z5121_assgn5121;
        z5121_assgn51211 <= z5121_assgn51210;
        z5121_assgn51212 <= z5121_assgn51211;
        z5121_assgn51213 <= z5121_assgn51212;
        z1811_assgn1811 <= z5121_assgn51213;
        z5151_assgn51510 <= z5151_assgn5151;
        z5151_assgn51511 <= z5151_assgn51510;
        z5151_assgn51512 <= z5151_assgn51511;
        z5151_assgn51513 <= z5151_assgn51512;
        z1839_assgn1839 <= z5151_assgn51513;
        z5155_assgn51550 <= z5155_assgn5155;
        z5155_assgn51551 <= z5155_assgn51550;
        z5155_assgn51552 <= z5155_assgn51551;
        z5155_assgn51553 <= z5155_assgn51552;
        z1841_assgn1841 <= z5155_assgn51553;
        z5163_assgn51630 <= z5163_assgn5163;
        z5163_assgn51631 <= z5163_assgn51630;
        z5163_assgn51632 <= z5163_assgn51631;
        z5163_assgn51633 <= z5163_assgn51632;
        z1847_assgn1847 <= z5163_assgn51633;
        z5167_assgn51670 <= z5167_assgn5167;
        z5167_assgn51671 <= z5167_assgn51670;
        z5167_assgn51672 <= z5167_assgn51671;
        z5167_assgn51673 <= z5167_assgn51672;
        z1849_assgn1849 <= z5167_assgn51673;
        u0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul1_G256_inv0;
        z5175_assgn51750 <= z5175_assgn5175;
        z5175_assgn51751 <= z5175_assgn51750;
        z5175_assgn51752 <= z5175_assgn51751;
        z5175_assgn51753 <= z5175_assgn51752;
        z1855_assgn1855 <= z5175_assgn51753;
        z5179_assgn51790 <= z5179_assgn5179;
        z5179_assgn51791 <= z5179_assgn51790;
        z5179_assgn51792 <= z5179_assgn51791;
        z5179_assgn51793 <= z5179_assgn51792;
        z1857_assgn1857 <= z5179_assgn51793;
        u1_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul1_G256_inv0;
        z5193_assgn51930 <= z5193_assgn5193;
        z5193_assgn51931 <= z5193_assgn51930;
        z5193_assgn51932 <= z5193_assgn51931;
        z5193_assgn51933 <= z5193_assgn51932;
        z1869_assgn1869 <= z5193_assgn51933;
        z5197_assgn51970 <= z5197_assgn5197;
        z5197_assgn51971 <= z5197_assgn51970;
        z5197_assgn51972 <= z5197_assgn51971;
        z5197_assgn51973 <= z5197_assgn51972;
        z1871_assgn1871 <= z5197_assgn51973;
        z5205_assgn52050 <= z5205_assgn5205;
        z5205_assgn52051 <= z5205_assgn52050;
        z5205_assgn52052 <= z5205_assgn52051;
        z5205_assgn52053 <= z5205_assgn52052;
        z1877_assgn1877 <= z5205_assgn52053;
        z5209_assgn52090 <= z5209_assgn5209;
        z5209_assgn52091 <= z5209_assgn52090;
        z5209_assgn52092 <= z5209_assgn52091;
        z5209_assgn52093 <= z5209_assgn52092;
        z1879_assgn1879 <= z5209_assgn52093;
        u0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul1_G256_inv0;
        z5217_assgn52170 <= z5217_assgn5217;
        z5217_assgn52171 <= z5217_assgn52170;
        z5217_assgn52172 <= z5217_assgn52171;
        z5217_assgn52173 <= z5217_assgn52172;
        z1885_assgn1885 <= z5217_assgn52173;
        z5221_assgn52210 <= z5221_assgn5221;
        z5221_assgn52211 <= z5221_assgn52210;
        z5221_assgn52212 <= z5221_assgn52211;
        z5221_assgn52213 <= z5221_assgn52212;
        z1887_assgn1887 <= z5221_assgn52213;
        u1_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul1_G256_inv0;
        z5239_assgn52390 <= z5239_assgn5239;
        z5239_assgn52391 <= z5239_assgn52390;
        z5239_assgn52392 <= z5239_assgn52391;
        z5239_assgn52393 <= z5239_assgn52392;
        z1903_assgn1903 <= z5239_assgn52393;
        z5243_assgn52430 <= z5243_assgn5243;
        z5243_assgn52431 <= z5243_assgn52430;
        z5243_assgn52432 <= z5243_assgn52431;
        z5243_assgn52433 <= z5243_assgn52432;
        z1905_assgn1905 <= z5243_assgn52433;
        z5251_assgn52510 <= z5251_assgn5251;
        z5251_assgn52511 <= z5251_assgn52510;
        z5251_assgn52512 <= z5251_assgn52511;
        z5251_assgn52513 <= z5251_assgn52512;
        z1911_assgn1911 <= z5251_assgn52513;
        z5255_assgn52550 <= z5255_assgn5255;
        z5255_assgn52551 <= z5255_assgn52550;
        z5255_assgn52552 <= z5255_assgn52551;
        z5255_assgn52553 <= z5255_assgn52552;
        z1913_assgn1913 <= z5255_assgn52553;
        u0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul1_G256_inv0;
        z5263_assgn52630 <= z5263_assgn5263;
        z5263_assgn52631 <= z5263_assgn52630;
        z5263_assgn52632 <= z5263_assgn52631;
        z5263_assgn52633 <= z5263_assgn52632;
        z1919_assgn1919 <= z5263_assgn52633;
        z5267_assgn52670 <= z5267_assgn5267;
        z5267_assgn52671 <= z5267_assgn52670;
        z5267_assgn52672 <= z5267_assgn52671;
        z5267_assgn52673 <= z5267_assgn52672;
        z1921_assgn1921 <= z5267_assgn52673;
        u1_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul1_G256_inv0;
        z5279_assgn52790 <= z5279_assgn5279;
        z5279_assgn52791 <= z5279_assgn52790;
        z5279_assgn52792 <= z5279_assgn52791;
        z5279_assgn52793 <= z5279_assgn52792;
        z5279_assgn52794 <= z5279_assgn52793;
        z1931_assgn1931 <= z5279_assgn52794;
        z5283_assgn52830 <= z5283_assgn5283;
        z5283_assgn52831 <= z5283_assgn52830;
        z5283_assgn52832 <= z5283_assgn52831;
        z5283_assgn52833 <= z5283_assgn52832;
        z5283_assgn52834 <= z5283_assgn52833;
        z1933_assgn1933 <= z5283_assgn52834;
        z5301_assgn53010 <= z5301_assgn5301;
        z5301_assgn53011 <= z5301_assgn53010;
        z5301_assgn53012 <= z5301_assgn53011;
        z5301_assgn53013 <= z5301_assgn53012;
        z1949_assgn1949 <= z5301_assgn53013;
        z5305_assgn53050 <= z5305_assgn5305;
        z5305_assgn53051 <= z5305_assgn53050;
        z5305_assgn53052 <= z5305_assgn53051;
        z5305_assgn53053 <= z5305_assgn53052;
        z1951_assgn1951 <= z5305_assgn53053;
        z5309_assgn53090 <= z5309_assgn5309;
        z5309_assgn53091 <= z5309_assgn53090;
        z5309_assgn53092 <= z5309_assgn53091;
        z5309_assgn53093 <= z5309_assgn53092;
        z1953_assgn1953 <= z5309_assgn53093;
        z5313_assgn53130 <= z5313_assgn5313;
        z5313_assgn53131 <= z5313_assgn53130;
        z5313_assgn53132 <= z5313_assgn53131;
        z5313_assgn53133 <= z5313_assgn53132;
        z1955_assgn1955 <= z5313_assgn53133;
        z5317_assgn53170 <= z5317_assgn5317;
        z5317_assgn53171 <= z5317_assgn53170;
        z5317_assgn53172 <= z5317_assgn53171;
        z5317_assgn53173 <= z5317_assgn53172;
        z1957_assgn1957 <= z5317_assgn53173;
        z5321_assgn53210 <= z5321_assgn5321;
        z5321_assgn53211 <= z5321_assgn53210;
        z5321_assgn53212 <= z5321_assgn53211;
        z5321_assgn53213 <= z5321_assgn53212;
        z1959_assgn1959 <= z5321_assgn53213;
        z5351_assgn53510 <= z5351_assgn5351;
        z5351_assgn53511 <= z5351_assgn53510;
        z5351_assgn53512 <= z5351_assgn53511;
        z5351_assgn53513 <= z5351_assgn53512;
        z1987_assgn1987 <= z5351_assgn53513;
        z5355_assgn53550 <= z5355_assgn5355;
        z5355_assgn53551 <= z5355_assgn53550;
        z5355_assgn53552 <= z5355_assgn53551;
        z5355_assgn53553 <= z5355_assgn53552;
        z1989_assgn1989 <= z5355_assgn53553;
        z5363_assgn53630 <= z5363_assgn5363;
        z5363_assgn53631 <= z5363_assgn53630;
        z5363_assgn53632 <= z5363_assgn53631;
        z5363_assgn53633 <= z5363_assgn53632;
        z1995_assgn1995 <= z5363_assgn53633;
        z5367_assgn53670 <= z5367_assgn5367;
        z5367_assgn53671 <= z5367_assgn53670;
        z5367_assgn53672 <= z5367_assgn53671;
        z5367_assgn53673 <= z5367_assgn53672;
        z1997_assgn1997 <= z5367_assgn53673;
        u0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul1_G256_inv0;
        z5375_assgn53750 <= z5375_assgn5375;
        z5375_assgn53751 <= z5375_assgn53750;
        z5375_assgn53752 <= z5375_assgn53751;
        z5375_assgn53753 <= z5375_assgn53752;
        z2003_assgn2003 <= z5375_assgn53753;
        z5379_assgn53790 <= z5379_assgn5379;
        z5379_assgn53791 <= z5379_assgn53790;
        z5379_assgn53792 <= z5379_assgn53791;
        z5379_assgn53793 <= z5379_assgn53792;
        z2005_assgn2005 <= z5379_assgn53793;
        u1_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul1_G256_inv0;
        z5393_assgn53930 <= z5393_assgn5393;
        z5393_assgn53931 <= z5393_assgn53930;
        z5393_assgn53932 <= z5393_assgn53931;
        z5393_assgn53933 <= z5393_assgn53932;
        z2017_assgn2017 <= z5393_assgn53933;
        z5397_assgn53970 <= z5397_assgn5397;
        z5397_assgn53971 <= z5397_assgn53970;
        z5397_assgn53972 <= z5397_assgn53971;
        z5397_assgn53973 <= z5397_assgn53972;
        z2019_assgn2019 <= z5397_assgn53973;
        z5405_assgn54050 <= z5405_assgn5405;
        z5405_assgn54051 <= z5405_assgn54050;
        z5405_assgn54052 <= z5405_assgn54051;
        z5405_assgn54053 <= z5405_assgn54052;
        z2025_assgn2025 <= z5405_assgn54053;
        z5409_assgn54090 <= z5409_assgn5409;
        z5409_assgn54091 <= z5409_assgn54090;
        z5409_assgn54092 <= z5409_assgn54091;
        z5409_assgn54093 <= z5409_assgn54092;
        z2027_assgn2027 <= z5409_assgn54093;
        u0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul1_G256_inv0;
        z5417_assgn54170 <= z5417_assgn5417;
        z5417_assgn54171 <= z5417_assgn54170;
        z5417_assgn54172 <= z5417_assgn54171;
        z5417_assgn54173 <= z5417_assgn54172;
        z2033_assgn2033 <= z5417_assgn54173;
        z5421_assgn54210 <= z5421_assgn5421;
        z5421_assgn54211 <= z5421_assgn54210;
        z5421_assgn54212 <= z5421_assgn54211;
        z5421_assgn54213 <= z5421_assgn54212;
        z2035_assgn2035 <= z5421_assgn54213;
        u1_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul1_G256_inv0;
        z5439_assgn54390 <= z5439_assgn5439;
        z5439_assgn54391 <= z5439_assgn54390;
        z5439_assgn54392 <= z5439_assgn54391;
        z5439_assgn54393 <= z5439_assgn54392;
        z2051_assgn2051 <= z5439_assgn54393;
        z5443_assgn54430 <= z5443_assgn5443;
        z5443_assgn54431 <= z5443_assgn54430;
        z5443_assgn54432 <= z5443_assgn54431;
        z5443_assgn54433 <= z5443_assgn54432;
        z2053_assgn2053 <= z5443_assgn54433;
        z5451_assgn54510 <= z5451_assgn5451;
        z5451_assgn54511 <= z5451_assgn54510;
        z5451_assgn54512 <= z5451_assgn54511;
        z5451_assgn54513 <= z5451_assgn54512;
        z2059_assgn2059 <= z5451_assgn54513;
        z5455_assgn54550 <= z5455_assgn5455;
        z5455_assgn54551 <= z5455_assgn54550;
        z5455_assgn54552 <= z5455_assgn54551;
        z5455_assgn54553 <= z5455_assgn54552;
        z2061_assgn2061 <= z5455_assgn54553;
        u0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul1_G256_inv0;
        z5463_assgn54630 <= z5463_assgn5463;
        z5463_assgn54631 <= z5463_assgn54630;
        z5463_assgn54632 <= z5463_assgn54631;
        z5463_assgn54633 <= z5463_assgn54632;
        z2067_assgn2067 <= z5463_assgn54633;
        z5467_assgn54670 <= z5467_assgn5467;
        z5467_assgn54671 <= z5467_assgn54670;
        z5467_assgn54672 <= z5467_assgn54671;
        z5467_assgn54673 <= z5467_assgn54672;
        z2069_assgn2069 <= z5467_assgn54673;
        u1_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul1_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul1_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul1_G256_inv0;
        z5479_assgn54790 <= z5479_assgn5479;
        z5479_assgn54791 <= z5479_assgn54790;
        z5479_assgn54792 <= z5479_assgn54791;
        z5479_assgn54793 <= z5479_assgn54792;
        z5479_assgn54794 <= z5479_assgn54793;
        z2079_assgn2079 <= z5479_assgn54794;
        z5483_assgn54830 <= z5483_assgn5483;
        z5483_assgn54831 <= z5483_assgn54830;
        z5483_assgn54832 <= z5483_assgn54831;
        z5483_assgn54833 <= z5483_assgn54832;
        z5483_assgn54834 <= z5483_assgn54833;
        z2081_assgn2081 <= z5483_assgn54834;
        z5495_assgn54950 <= z5495_assgn5495;
        z5495_assgn54951 <= z5495_assgn54950;
        z5495_assgn54952 <= z5495_assgn54951;
        z5495_assgn54953 <= z5495_assgn54952;
        z5495_assgn54954 <= z5495_assgn54953;
        z2091_assgn2091 <= z5495_assgn54954;
        z5499_assgn54990 <= z5499_assgn5499;
        z5499_assgn54991 <= z5499_assgn54990;
        z5499_assgn54992 <= z5499_assgn54991;
        z5499_assgn54993 <= z5499_assgn54992;
        z5499_assgn54994 <= z5499_assgn54993;
        z2093_assgn2093 <= z5499_assgn54994;
        z5525_assgn55250 <= z5525_assgn5525;
        z5525_assgn55251 <= z5525_assgn55250;
        z5525_assgn55252 <= z5525_assgn55251;
        z5525_assgn55253 <= z5525_assgn55252;
        z2117_assgn2117 <= z5525_assgn55253;
        z5529_assgn55290 <= z5529_assgn5529;
        z5529_assgn55291 <= z5529_assgn55290;
        z5529_assgn55292 <= z5529_assgn55291;
        z5529_assgn55293 <= z5529_assgn55292;
        z2119_assgn2119 <= z5529_assgn55293;
        z5533_assgn55330 <= z5533_assgn5533;
        z5533_assgn55331 <= z5533_assgn55330;
        z5533_assgn55332 <= z5533_assgn55331;
        z5533_assgn55333 <= z5533_assgn55332;
        z2121_assgn2121 <= z5533_assgn55333;
        z5537_assgn55370 <= z5537_assgn5537;
        z5537_assgn55371 <= z5537_assgn55370;
        z5537_assgn55372 <= z5537_assgn55371;
        z5537_assgn55373 <= z5537_assgn55372;
        z2123_assgn2123 <= z5537_assgn55373;
        z5541_assgn55410 <= z5541_assgn5541;
        z5541_assgn55411 <= z5541_assgn55410;
        z5541_assgn55412 <= z5541_assgn55411;
        z5541_assgn55413 <= z5541_assgn55412;
        z2125_assgn2125 <= z5541_assgn55413;
        z5545_assgn55450 <= z5545_assgn5545;
        z5545_assgn55451 <= z5545_assgn55450;
        z5545_assgn55452 <= z5545_assgn55451;
        z5545_assgn55453 <= z5545_assgn55452;
        z2127_assgn2127 <= z5545_assgn55453;
        z5575_assgn55750 <= z5575_assgn5575;
        z5575_assgn55751 <= z5575_assgn55750;
        z5575_assgn55752 <= z5575_assgn55751;
        z5575_assgn55753 <= z5575_assgn55752;
        z2155_assgn2155 <= z5575_assgn55753;
        z5579_assgn55790 <= z5579_assgn5579;
        z5579_assgn55791 <= z5579_assgn55790;
        z5579_assgn55792 <= z5579_assgn55791;
        z5579_assgn55793 <= z5579_assgn55792;
        z2157_assgn2157 <= z5579_assgn55793;
        z5583_assgn55830 <= z5583_assgn5583;
        z5583_assgn55831 <= z5583_assgn55830;
        z5583_assgn55832 <= z5583_assgn55831;
        z5583_assgn55833 <= z5583_assgn55832;
        z2159_assgn2159 <= z5583_assgn55833;
        z5587_assgn55870 <= z5587_assgn5587;
        z5587_assgn55871 <= z5587_assgn55870;
        z5587_assgn55872 <= z5587_assgn55871;
        z5587_assgn55873 <= z5587_assgn55872;
        z2161_assgn2161 <= z5587_assgn55873;
        z5591_assgn55910 <= z5591_assgn5591;
        z5591_assgn55911 <= z5591_assgn55910;
        z5591_assgn55912 <= z5591_assgn55911;
        z5591_assgn55913 <= z5591_assgn55912;
        z2163_assgn2163 <= z5591_assgn55913;
        z5595_assgn55950 <= z5595_assgn5595;
        z5595_assgn55951 <= z5595_assgn55950;
        z5595_assgn55952 <= z5595_assgn55951;
        z5595_assgn55953 <= z5595_assgn55952;
        z2165_assgn2165 <= z5595_assgn55953;
        z5625_assgn56250 <= z5625_assgn5625;
        z5625_assgn56251 <= z5625_assgn56250;
        z5625_assgn56252 <= z5625_assgn56251;
        z5625_assgn56253 <= z5625_assgn56252;
        z2193_assgn2193 <= z5625_assgn56253;
        z5629_assgn56290 <= z5629_assgn5629;
        z5629_assgn56291 <= z5629_assgn56290;
        z5629_assgn56292 <= z5629_assgn56291;
        z5629_assgn56293 <= z5629_assgn56292;
        z2195_assgn2195 <= z5629_assgn56293;
        z5637_assgn56370 <= z5637_assgn5637;
        z5637_assgn56371 <= z5637_assgn56370;
        z5637_assgn56372 <= z5637_assgn56371;
        z5637_assgn56373 <= z5637_assgn56372;
        z2201_assgn2201 <= z5637_assgn56373;
        z5641_assgn56410 <= z5641_assgn5641;
        z5641_assgn56411 <= z5641_assgn56410;
        z5641_assgn56412 <= z5641_assgn56411;
        z5641_assgn56413 <= z5641_assgn56412;
        z2203_assgn2203 <= z5641_assgn56413;
        u0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul0_G16_mul2_G256_inv0;
        z5649_assgn56490 <= z5649_assgn5649;
        z5649_assgn56491 <= z5649_assgn56490;
        z5649_assgn56492 <= z5649_assgn56491;
        z5649_assgn56493 <= z5649_assgn56492;
        z2209_assgn2209 <= z5649_assgn56493;
        z5653_assgn56530 <= z5653_assgn5653;
        z5653_assgn56531 <= z5653_assgn56530;
        z5653_assgn56532 <= z5653_assgn56531;
        z5653_assgn56533 <= z5653_assgn56532;
        z2211_assgn2211 <= z5653_assgn56533;
        u1_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul0_G16_mul2_G256_inv0;
        z5667_assgn56670 <= z5667_assgn5667;
        z5667_assgn56671 <= z5667_assgn56670;
        z5667_assgn56672 <= z5667_assgn56671;
        z5667_assgn56673 <= z5667_assgn56672;
        z2223_assgn2223 <= z5667_assgn56673;
        z5671_assgn56710 <= z5671_assgn5671;
        z5671_assgn56711 <= z5671_assgn56710;
        z5671_assgn56712 <= z5671_assgn56711;
        z5671_assgn56713 <= z5671_assgn56712;
        z2225_assgn2225 <= z5671_assgn56713;
        z5679_assgn56790 <= z5679_assgn5679;
        z5679_assgn56791 <= z5679_assgn56790;
        z5679_assgn56792 <= z5679_assgn56791;
        z5679_assgn56793 <= z5679_assgn56792;
        z2231_assgn2231 <= z5679_assgn56793;
        z5683_assgn56830 <= z5683_assgn5683;
        z5683_assgn56831 <= z5683_assgn56830;
        z5683_assgn56832 <= z5683_assgn56831;
        z5683_assgn56833 <= z5683_assgn56832;
        z2233_assgn2233 <= z5683_assgn56833;
        u0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul0_G16_mul2_G256_inv0;
        z5691_assgn56910 <= z5691_assgn5691;
        z5691_assgn56911 <= z5691_assgn56910;
        z5691_assgn56912 <= z5691_assgn56911;
        z5691_assgn56913 <= z5691_assgn56912;
        z2239_assgn2239 <= z5691_assgn56913;
        z5695_assgn56950 <= z5695_assgn5695;
        z5695_assgn56951 <= z5695_assgn56950;
        z5695_assgn56952 <= z5695_assgn56951;
        z5695_assgn56953 <= z5695_assgn56952;
        z2241_assgn2241 <= z5695_assgn56953;
        u1_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul0_G16_mul2_G256_inv0;
        z5713_assgn57130 <= z5713_assgn5713;
        z5713_assgn57131 <= z5713_assgn57130;
        z5713_assgn57132 <= z5713_assgn57131;
        z5713_assgn57133 <= z5713_assgn57132;
        z2257_assgn2257 <= z5713_assgn57133;
        z5717_assgn57170 <= z5717_assgn5717;
        z5717_assgn57171 <= z5717_assgn57170;
        z5717_assgn57172 <= z5717_assgn57171;
        z5717_assgn57173 <= z5717_assgn57172;
        z2259_assgn2259 <= z5717_assgn57173;
        z5725_assgn57250 <= z5725_assgn5725;
        z5725_assgn57251 <= z5725_assgn57250;
        z5725_assgn57252 <= z5725_assgn57251;
        z5725_assgn57253 <= z5725_assgn57252;
        z2265_assgn2265 <= z5725_assgn57253;
        z5729_assgn57290 <= z5729_assgn5729;
        z5729_assgn57291 <= z5729_assgn57290;
        z5729_assgn57292 <= z5729_assgn57291;
        z5729_assgn57293 <= z5729_assgn57292;
        z2267_assgn2267 <= z5729_assgn57293;
        u0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul0_G16_mul2_G256_inv0;
        z5737_assgn57370 <= z5737_assgn5737;
        z5737_assgn57371 <= z5737_assgn57370;
        z5737_assgn57372 <= z5737_assgn57371;
        z5737_assgn57373 <= z5737_assgn57372;
        z2273_assgn2273 <= z5737_assgn57373;
        z5741_assgn57410 <= z5741_assgn5741;
        z5741_assgn57411 <= z5741_assgn57410;
        z5741_assgn57412 <= z5741_assgn57411;
        z5741_assgn57413 <= z5741_assgn57412;
        z2275_assgn2275 <= z5741_assgn57413;
        u1_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul0_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul0_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul0_G16_mul2_G256_inv0;
        z5753_assgn57530 <= z5753_assgn5753;
        z5753_assgn57531 <= z5753_assgn57530;
        z5753_assgn57532 <= z5753_assgn57531;
        z5753_assgn57533 <= z5753_assgn57532;
        z5753_assgn57534 <= z5753_assgn57533;
        z2285_assgn2285 <= z5753_assgn57534;
        z5757_assgn57570 <= z5757_assgn5757;
        z5757_assgn57571 <= z5757_assgn57570;
        z5757_assgn57572 <= z5757_assgn57571;
        z5757_assgn57573 <= z5757_assgn57572;
        z5757_assgn57574 <= z5757_assgn57573;
        z2287_assgn2287 <= z5757_assgn57574;
        z5765_assgn57650 <= z5765_assgn5765;
        z5765_assgn57651 <= z5765_assgn57650;
        z5765_assgn57652 <= z5765_assgn57651;
        z5765_assgn57653 <= z5765_assgn57652;
        z5765_assgn57654 <= z5765_assgn57653;
        z2293_assgn2293 <= z5765_assgn57654;
        z5769_assgn57690 <= z5769_assgn5769;
        z5769_assgn57691 <= z5769_assgn57690;
        z5769_assgn57692 <= z5769_assgn57691;
        z5769_assgn57693 <= z5769_assgn57692;
        z5769_assgn57694 <= z5769_assgn57693;
        z2295_assgn2295 <= z5769_assgn57694;
        z5773_assgn57730 <= z5773_assgn5773;
        z5773_assgn57731 <= z5773_assgn57730;
        z5773_assgn57732 <= z5773_assgn57731;
        z5773_assgn57733 <= z5773_assgn57732;
        z5773_assgn57734 <= z5773_assgn57733;
        z2297_assgn2297 <= z5773_assgn57734;
        z5777_assgn57770 <= z5777_assgn5777;
        z5777_assgn57771 <= z5777_assgn57770;
        z5777_assgn57772 <= z5777_assgn57771;
        z5777_assgn57773 <= z5777_assgn57772;
        z5777_assgn57774 <= z5777_assgn57773;
        z2299_assgn2299 <= z5777_assgn57774;
        z5781_assgn57810 <= z5781_assgn5781;
        z5781_assgn57811 <= z5781_assgn57810;
        z5781_assgn57812 <= z5781_assgn57811;
        z5781_assgn57813 <= z5781_assgn57812;
        z5781_assgn57814 <= z5781_assgn57813;
        z2301_assgn2301 <= z5781_assgn57814;
        z5785_assgn57850 <= z5785_assgn5785;
        z5785_assgn57851 <= z5785_assgn57850;
        z5785_assgn57852 <= z5785_assgn57851;
        z5785_assgn57853 <= z5785_assgn57852;
        z5785_assgn57854 <= z5785_assgn57853;
        z2303_assgn2303 <= z5785_assgn57854;
        z5797_assgn57970 <= z5797_assgn5797;
        z5797_assgn57971 <= z5797_assgn57970;
        z5797_assgn57972 <= z5797_assgn57971;
        z5797_assgn57973 <= z5797_assgn57972;
        z5797_assgn57974 <= z5797_assgn57973;
        z2313_assgn2313 <= z5797_assgn57974;
        z5801_assgn58010 <= z5801_assgn5801;
        z5801_assgn58011 <= z5801_assgn58010;
        z5801_assgn58012 <= z5801_assgn58011;
        z5801_assgn58013 <= z5801_assgn58012;
        z5801_assgn58014 <= z5801_assgn58013;
        z2315_assgn2315 <= z5801_assgn58014;
        z5815_assgn58150 <= z5815_assgn5815;
        z5815_assgn58151 <= z5815_assgn58150;
        z5815_assgn58152 <= z5815_assgn58151;
        z5815_assgn58153 <= z5815_assgn58152;
        z2327_assgn2327 <= z5815_assgn58153;
        z5819_assgn58190 <= z5819_assgn5819;
        z5819_assgn58191 <= z5819_assgn58190;
        z5819_assgn58192 <= z5819_assgn58191;
        z5819_assgn58193 <= z5819_assgn58192;
        z2329_assgn2329 <= z5819_assgn58193;
        z5823_assgn58230 <= z5823_assgn5823;
        z5823_assgn58231 <= z5823_assgn58230;
        z5823_assgn58232 <= z5823_assgn58231;
        z5823_assgn58233 <= z5823_assgn58232;
        z2331_assgn2331 <= z5823_assgn58233;
        z5827_assgn58270 <= z5827_assgn5827;
        z5827_assgn58271 <= z5827_assgn58270;
        z5827_assgn58272 <= z5827_assgn58271;
        z5827_assgn58273 <= z5827_assgn58272;
        z2333_assgn2333 <= z5827_assgn58273;
        z5831_assgn58310 <= z5831_assgn5831;
        z5831_assgn58311 <= z5831_assgn58310;
        z5831_assgn58312 <= z5831_assgn58311;
        z5831_assgn58313 <= z5831_assgn58312;
        z2335_assgn2335 <= z5831_assgn58313;
        z5835_assgn58350 <= z5835_assgn5835;
        z5835_assgn58351 <= z5835_assgn58350;
        z5835_assgn58352 <= z5835_assgn58351;
        z5835_assgn58353 <= z5835_assgn58352;
        z2337_assgn2337 <= z5835_assgn58353;
        z5865_assgn58650 <= z5865_assgn5865;
        z5865_assgn58651 <= z5865_assgn58650;
        z5865_assgn58652 <= z5865_assgn58651;
        z5865_assgn58653 <= z5865_assgn58652;
        z2365_assgn2365 <= z5865_assgn58653;
        z5869_assgn58690 <= z5869_assgn5869;
        z5869_assgn58691 <= z5869_assgn58690;
        z5869_assgn58692 <= z5869_assgn58691;
        z5869_assgn58693 <= z5869_assgn58692;
        z2367_assgn2367 <= z5869_assgn58693;
        z5877_assgn58770 <= z5877_assgn5877;
        z5877_assgn58771 <= z5877_assgn58770;
        z5877_assgn58772 <= z5877_assgn58771;
        z5877_assgn58773 <= z5877_assgn58772;
        z2373_assgn2373 <= z5877_assgn58773;
        z5881_assgn58810 <= z5881_assgn5881;
        z5881_assgn58811 <= z5881_assgn58810;
        z5881_assgn58812 <= z5881_assgn58811;
        z5881_assgn58813 <= z5881_assgn58812;
        z2375_assgn2375 <= z5881_assgn58813;
        u0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul1_G16_mul2_G256_inv0;
        z5889_assgn58890 <= z5889_assgn5889;
        z5889_assgn58891 <= z5889_assgn58890;
        z5889_assgn58892 <= z5889_assgn58891;
        z5889_assgn58893 <= z5889_assgn58892;
        z2381_assgn2381 <= z5889_assgn58893;
        z5893_assgn58930 <= z5893_assgn5893;
        z5893_assgn58931 <= z5893_assgn58930;
        z5893_assgn58932 <= z5893_assgn58931;
        z5893_assgn58933 <= z5893_assgn58932;
        z2383_assgn2383 <= z5893_assgn58933;
        u1_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul1_G16_mul2_G256_inv0;
        z5907_assgn59070 <= z5907_assgn5907;
        z5907_assgn59071 <= z5907_assgn59070;
        z5907_assgn59072 <= z5907_assgn59071;
        z5907_assgn59073 <= z5907_assgn59072;
        z2395_assgn2395 <= z5907_assgn59073;
        z5911_assgn59110 <= z5911_assgn5911;
        z5911_assgn59111 <= z5911_assgn59110;
        z5911_assgn59112 <= z5911_assgn59111;
        z5911_assgn59113 <= z5911_assgn59112;
        z2397_assgn2397 <= z5911_assgn59113;
        z5919_assgn59190 <= z5919_assgn5919;
        z5919_assgn59191 <= z5919_assgn59190;
        z5919_assgn59192 <= z5919_assgn59191;
        z5919_assgn59193 <= z5919_assgn59192;
        z2403_assgn2403 <= z5919_assgn59193;
        z5923_assgn59230 <= z5923_assgn5923;
        z5923_assgn59231 <= z5923_assgn59230;
        z5923_assgn59232 <= z5923_assgn59231;
        z5923_assgn59233 <= z5923_assgn59232;
        z2405_assgn2405 <= z5923_assgn59233;
        u0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul1_G16_mul2_G256_inv0;
        z5931_assgn59310 <= z5931_assgn5931;
        z5931_assgn59311 <= z5931_assgn59310;
        z5931_assgn59312 <= z5931_assgn59311;
        z5931_assgn59313 <= z5931_assgn59312;
        z2411_assgn2411 <= z5931_assgn59313;
        z5935_assgn59350 <= z5935_assgn5935;
        z5935_assgn59351 <= z5935_assgn59350;
        z5935_assgn59352 <= z5935_assgn59351;
        z5935_assgn59353 <= z5935_assgn59352;
        z2413_assgn2413 <= z5935_assgn59353;
        u1_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul1_G16_mul2_G256_inv0;
        z5953_assgn59530 <= z5953_assgn5953;
        z5953_assgn59531 <= z5953_assgn59530;
        z5953_assgn59532 <= z5953_assgn59531;
        z5953_assgn59533 <= z5953_assgn59532;
        z2429_assgn2429 <= z5953_assgn59533;
        z5957_assgn59570 <= z5957_assgn5957;
        z5957_assgn59571 <= z5957_assgn59570;
        z5957_assgn59572 <= z5957_assgn59571;
        z5957_assgn59573 <= z5957_assgn59572;
        z2431_assgn2431 <= z5957_assgn59573;
        z5965_assgn59650 <= z5965_assgn5965;
        z5965_assgn59651 <= z5965_assgn59650;
        z5965_assgn59652 <= z5965_assgn59651;
        z5965_assgn59653 <= z5965_assgn59652;
        z2437_assgn2437 <= z5965_assgn59653;
        z5969_assgn59690 <= z5969_assgn5969;
        z5969_assgn59691 <= z5969_assgn59690;
        z5969_assgn59692 <= z5969_assgn59691;
        z5969_assgn59693 <= z5969_assgn59692;
        z2439_assgn2439 <= z5969_assgn59693;
        u0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul1_G16_mul2_G256_inv0;
        z5977_assgn59770 <= z5977_assgn5977;
        z5977_assgn59771 <= z5977_assgn59770;
        z5977_assgn59772 <= z5977_assgn59771;
        z5977_assgn59773 <= z5977_assgn59772;
        z2445_assgn2445 <= z5977_assgn59773;
        z5981_assgn59810 <= z5981_assgn5981;
        z5981_assgn59811 <= z5981_assgn59810;
        z5981_assgn59812 <= z5981_assgn59811;
        z5981_assgn59813 <= z5981_assgn59812;
        z2447_assgn2447 <= z5981_assgn59813;
        u1_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul1_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul1_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul1_G16_mul2_G256_inv0;
        z5993_assgn59930 <= z5993_assgn5993;
        z5993_assgn59931 <= z5993_assgn59930;
        z5993_assgn59932 <= z5993_assgn59931;
        z5993_assgn59933 <= z5993_assgn59932;
        z5993_assgn59934 <= z5993_assgn59933;
        z2457_assgn2457 <= z5993_assgn59934;
        z5997_assgn59970 <= z5997_assgn5997;
        z5997_assgn59971 <= z5997_assgn59970;
        z5997_assgn59972 <= z5997_assgn59971;
        z5997_assgn59973 <= z5997_assgn59972;
        z5997_assgn59974 <= z5997_assgn59973;
        z2459_assgn2459 <= z5997_assgn59974;
        z6015_assgn60150 <= z6015_assgn6015;
        z6015_assgn60151 <= z6015_assgn60150;
        z6015_assgn60152 <= z6015_assgn60151;
        z6015_assgn60153 <= z6015_assgn60152;
        z2475_assgn2475 <= z6015_assgn60153;
        z6019_assgn60190 <= z6019_assgn6019;
        z6019_assgn60191 <= z6019_assgn60190;
        z6019_assgn60192 <= z6019_assgn60191;
        z6019_assgn60193 <= z6019_assgn60192;
        z2477_assgn2477 <= z6019_assgn60193;
        z6023_assgn60230 <= z6023_assgn6023;
        z6023_assgn60231 <= z6023_assgn60230;
        z6023_assgn60232 <= z6023_assgn60231;
        z6023_assgn60233 <= z6023_assgn60232;
        z2479_assgn2479 <= z6023_assgn60233;
        z6027_assgn60270 <= z6027_assgn6027;
        z6027_assgn60271 <= z6027_assgn60270;
        z6027_assgn60272 <= z6027_assgn60271;
        z6027_assgn60273 <= z6027_assgn60272;
        z2481_assgn2481 <= z6027_assgn60273;
        z6031_assgn60310 <= z6031_assgn6031;
        z6031_assgn60311 <= z6031_assgn60310;
        z6031_assgn60312 <= z6031_assgn60311;
        z6031_assgn60313 <= z6031_assgn60312;
        z2483_assgn2483 <= z6031_assgn60313;
        z6035_assgn60350 <= z6035_assgn6035;
        z6035_assgn60351 <= z6035_assgn60350;
        z6035_assgn60352 <= z6035_assgn60351;
        z6035_assgn60353 <= z6035_assgn60352;
        z2485_assgn2485 <= z6035_assgn60353;
        z6065_assgn60650 <= z6065_assgn6065;
        z6065_assgn60651 <= z6065_assgn60650;
        z6065_assgn60652 <= z6065_assgn60651;
        z6065_assgn60653 <= z6065_assgn60652;
        z2513_assgn2513 <= z6065_assgn60653;
        z6069_assgn60690 <= z6069_assgn6069;
        z6069_assgn60691 <= z6069_assgn60690;
        z6069_assgn60692 <= z6069_assgn60691;
        z6069_assgn60693 <= z6069_assgn60692;
        z2515_assgn2515 <= z6069_assgn60693;
        z6077_assgn60770 <= z6077_assgn6077;
        z6077_assgn60771 <= z6077_assgn60770;
        z6077_assgn60772 <= z6077_assgn60771;
        z6077_assgn60773 <= z6077_assgn60772;
        z2521_assgn2521 <= z6077_assgn60773;
        z6081_assgn60810 <= z6081_assgn6081;
        z6081_assgn60811 <= z6081_assgn60810;
        z6081_assgn60812 <= z6081_assgn60811;
        z6081_assgn60813 <= z6081_assgn60812;
        z2523_assgn2523 <= z6081_assgn60813;
        u0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc20_G4_mul2_G16_mul2_G256_inv0;
        z6089_assgn60890 <= z6089_assgn6089;
        z6089_assgn60891 <= z6089_assgn60890;
        z6089_assgn60892 <= z6089_assgn60891;
        z6089_assgn60893 <= z6089_assgn60892;
        z2529_assgn2529 <= z6089_assgn60893;
        z6093_assgn60930 <= z6093_assgn6093;
        z6093_assgn60931 <= z6093_assgn60930;
        z6093_assgn60932 <= z6093_assgn60931;
        z6093_assgn60933 <= z6093_assgn60932;
        z2531_assgn2531 <= z6093_assgn60933;
        u1_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc20_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc20_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc20_G4_mul2_G16_mul2_G256_inv0;
        z6107_assgn61070 <= z6107_assgn6107;
        z6107_assgn61071 <= z6107_assgn61070;
        z6107_assgn61072 <= z6107_assgn61071;
        z6107_assgn61073 <= z6107_assgn61072;
        z2543_assgn2543 <= z6107_assgn61073;
        z6111_assgn61110 <= z6111_assgn6111;
        z6111_assgn61111 <= z6111_assgn61110;
        z6111_assgn61112 <= z6111_assgn61111;
        z6111_assgn61113 <= z6111_assgn61112;
        z2545_assgn2545 <= z6111_assgn61113;
        z6119_assgn61190 <= z6119_assgn6119;
        z6119_assgn61191 <= z6119_assgn61190;
        z6119_assgn61192 <= z6119_assgn61191;
        z6119_assgn61193 <= z6119_assgn61192;
        z2551_assgn2551 <= z6119_assgn61193;
        z6123_assgn61230 <= z6123_assgn6123;
        z6123_assgn61231 <= z6123_assgn61230;
        z6123_assgn61232 <= z6123_assgn61231;
        z6123_assgn61233 <= z6123_assgn61232;
        z2553_assgn2553 <= z6123_assgn61233;
        u0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc21_G4_mul2_G16_mul2_G256_inv0;
        z6131_assgn61310 <= z6131_assgn6131;
        z6131_assgn61311 <= z6131_assgn61310;
        z6131_assgn61312 <= z6131_assgn61311;
        z6131_assgn61313 <= z6131_assgn61312;
        z2559_assgn2559 <= z6131_assgn61313;
        z6135_assgn61350 <= z6135_assgn6135;
        z6135_assgn61351 <= z6135_assgn61350;
        z6135_assgn61352 <= z6135_assgn61351;
        z6135_assgn61353 <= z6135_assgn61352;
        z2561_assgn2561 <= z6135_assgn61353;
        u1_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc21_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc21_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc21_G4_mul2_G16_mul2_G256_inv0;
        z6153_assgn61530 <= z6153_assgn6153;
        z6153_assgn61531 <= z6153_assgn61530;
        z6153_assgn61532 <= z6153_assgn61531;
        z6153_assgn61533 <= z6153_assgn61532;
        z2577_assgn2577 <= z6153_assgn61533;
        z6157_assgn61570 <= z6157_assgn6157;
        z6157_assgn61571 <= z6157_assgn61570;
        z6157_assgn61572 <= z6157_assgn61571;
        z6157_assgn61573 <= z6157_assgn61572;
        z2579_assgn2579 <= z6157_assgn61573;
        z6165_assgn61650 <= z6165_assgn6165;
        z6165_assgn61651 <= z6165_assgn61650;
        z6165_assgn61652 <= z6165_assgn61651;
        z6165_assgn61653 <= z6165_assgn61652;
        z2585_assgn2585 <= z6165_assgn61653;
        z6169_assgn61690 <= z6169_assgn6169;
        z6169_assgn61691 <= z6169_assgn61690;
        z6169_assgn61692 <= z6169_assgn61691;
        z6169_assgn61693 <= z6169_assgn61692;
        z2587_assgn2587 <= z6169_assgn61693;
        u0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= u0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p1_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p0_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p0_hpc22_G4_mul2_G16_mul2_G256_inv0;
        z6177_assgn61770 <= z6177_assgn6177;
        z6177_assgn61771 <= z6177_assgn61770;
        z6177_assgn61772 <= z6177_assgn61771;
        z6177_assgn61773 <= z6177_assgn61772;
        z2593_assgn2593 <= z6177_assgn61773;
        z6181_assgn61810 <= z6181_assgn6181;
        z6181_assgn61811 <= z6181_assgn61810;
        z6181_assgn61812 <= z6181_assgn61811;
        z6181_assgn61813 <= z6181_assgn61812;
        z2595_assgn2595 <= z6181_assgn61813;
        u1_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= u1_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p3_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p3_hpc22_G4_mul2_G16_mul2_G256_inv0;
        p2_hpc22_G4_mul2_G16_mul2_G256_inv0_reg <= p2_hpc22_G4_mul2_G16_mul2_G256_inv0;
        z6193_assgn61930 <= z6193_assgn6193;
        z6193_assgn61931 <= z6193_assgn61930;
        z6193_assgn61932 <= z6193_assgn61931;
        z6193_assgn61933 <= z6193_assgn61932;
        z6193_assgn61934 <= z6193_assgn61933;
        z2605_assgn2605 <= z6193_assgn61934;
        z6197_assgn61970 <= z6197_assgn6197;
        z6197_assgn61971 <= z6197_assgn61970;
        z6197_assgn61972 <= z6197_assgn61971;
        z6197_assgn61973 <= z6197_assgn61972;
        z6197_assgn61974 <= z6197_assgn61973;
        z2607_assgn2607 <= z6197_assgn61974;
        z6209_assgn62090 <= z6209_assgn6209;
        z6209_assgn62091 <= z6209_assgn62090;
        z6209_assgn62092 <= z6209_assgn62091;
        z6209_assgn62093 <= z6209_assgn62092;
        z6209_assgn62094 <= z6209_assgn62093;
        z2617_assgn2617 <= z6209_assgn62094;
        z6213_assgn62130 <= z6213_assgn6213;
        z6213_assgn62131 <= z6213_assgn62130;
        z6213_assgn62132 <= z6213_assgn62131;
        z6213_assgn62133 <= z6213_assgn62132;
        z6213_assgn62134 <= z6213_assgn62133;
        z2619_assgn2619 <= z6213_assgn62134;
        z6221_assgn62210 <= z6221_assgn6221;
        z6221_assgn62211 <= z6221_assgn62210;
        z6221_assgn62212 <= z6221_assgn62211;
        z6221_assgn62213 <= z6221_assgn62212;
        z6221_assgn62214 <= z6221_assgn62213;
        z2625_assgn2625 <= z6221_assgn62214;
        z6225_assgn62250 <= z6225_assgn6225;
        z6225_assgn62251 <= z6225_assgn62250;
        z6225_assgn62252 <= z6225_assgn62251;
        z6225_assgn62253 <= z6225_assgn62252;
        z6225_assgn62254 <= z6225_assgn62253;
        z2627_assgn2627 <= z6225_assgn62254;
        z6237_assgn62370 <= z6237_assgn6237;
        z6237_assgn62371 <= z6237_assgn62370;
        z6237_assgn62372 <= z6237_assgn62371;
        z6237_assgn62373 <= z6237_assgn62372;
        z6237_assgn62374 <= z6237_assgn62373;
        z2637_assgn2637 <= z6237_assgn62374;
        z6245_assgn62450 <= z6245_assgn6245;
        z6245_assgn62451 <= z6245_assgn62450;
        z6245_assgn62452 <= z6245_assgn62451;
        z6245_assgn62453 <= z6245_assgn62452;
        z6245_assgn62454 <= z6245_assgn62453;
        z2643_assgn2643 <= z6245_assgn62454;
        z6249_assgn62490 <= z6249_assgn6249;
        z6249_assgn62491 <= z6249_assgn62490;
        z6249_assgn62492 <= z6249_assgn62491;
        z6249_assgn62493 <= z6249_assgn62492;
        z6249_assgn62494 <= z6249_assgn62493;
        z2646_assgn2646 <= z6249_assgn62494;
        z6255_assgn62550 <= z6255_assgn6255;
        z6255_assgn62551 <= z6255_assgn62550;
        z6255_assgn62552 <= z6255_assgn62551;
        z6255_assgn62553 <= z6255_assgn62552;
        z6255_assgn62554 <= z6255_assgn62553;
        z2649_assgn2649 <= z6255_assgn62554;
        z6261_assgn62610 <= z6261_assgn6261;
        z6261_assgn62611 <= z6261_assgn62610;
        z6261_assgn62612 <= z6261_assgn62611;
        z6261_assgn62613 <= z6261_assgn62612;
        z6261_assgn62614 <= z6261_assgn62613;
        z2653_assgn2653 <= z6261_assgn62614;
        z6267_assgn62670 <= z6267_assgn6267;
        z6267_assgn62671 <= z6267_assgn62670;
        z6267_assgn62672 <= z6267_assgn62671;
        z6267_assgn62673 <= z6267_assgn62672;
        z6267_assgn62674 <= z6267_assgn62673;
        z2657_assgn2657 <= z6267_assgn62674;
        z6277_assgn62770 <= z6277_assgn6277;
        z6277_assgn62771 <= z6277_assgn62770;
        z6277_assgn62772 <= z6277_assgn62771;
        z6277_assgn62773 <= z6277_assgn62772;
        z6277_assgn62774 <= z6277_assgn62773;
        z2665_assgn2665 <= z6277_assgn62774;
        z6283_assgn62830 <= z6283_assgn6283;
        z6283_assgn62831 <= z6283_assgn62830;
        z6283_assgn62832 <= z6283_assgn62831;
        z6283_assgn62833 <= z6283_assgn62832;
        z6283_assgn62834 <= z6283_assgn62833;
        z2669_assgn2669 <= z6283_assgn62834;
        z6289_assgn62890 <= z6289_assgn6289;
        z6289_assgn62891 <= z6289_assgn62890;
        z6289_assgn62892 <= z6289_assgn62891;
        z6289_assgn62893 <= z6289_assgn62892;
        z6289_assgn62894 <= z6289_assgn62893;
        z2673_assgn2673 <= z6289_assgn62894;
        z6299_assgn62990 <= z6299_assgn6299;
        z6299_assgn62991 <= z6299_assgn62990;
        z6299_assgn62992 <= z6299_assgn62991;
        z6299_assgn62993 <= z6299_assgn62992;
        z6299_assgn62994 <= z6299_assgn62993;
        z2681_assgn2681 <= z6299_assgn62994;
        z6305_assgn63050 <= z6305_assgn6305;
        z6305_assgn63051 <= z6305_assgn63050;
        z6305_assgn63052 <= z6305_assgn63051;
        z6305_assgn63053 <= z6305_assgn63052;
        z6305_assgn63054 <= z6305_assgn63053;
        z2685_assgn2685 <= z6305_assgn63054;
        z6311_assgn63110 <= z6311_assgn6311;
        z6311_assgn63111 <= z6311_assgn63110;
        z6311_assgn63112 <= z6311_assgn63111;
        z6311_assgn63113 <= z6311_assgn63112;
        z6311_assgn63114 <= z6311_assgn63113;
        z2689_assgn2689 <= z6311_assgn63114;
        z6321_assgn63210 <= z6321_assgn6321;
        z6321_assgn63211 <= z6321_assgn63210;
        z6321_assgn63212 <= z6321_assgn63211;
        z6321_assgn63213 <= z6321_assgn63212;
        z6321_assgn63214 <= z6321_assgn63213;
        z2697_assgn2697 <= z6321_assgn63214;
        z6327_assgn63270 <= z6327_assgn6327;
        z6327_assgn63271 <= z6327_assgn63270;
        z6327_assgn63272 <= z6327_assgn63271;
        z6327_assgn63273 <= z6327_assgn63272;
        z6327_assgn63274 <= z6327_assgn63273;
        z2701_assgn2701 <= z6327_assgn63274;
        z6333_assgn63330 <= z6333_assgn6333;
        z6333_assgn63331 <= z6333_assgn63330;
        z6333_assgn63332 <= z6333_assgn63331;
        z6333_assgn63333 <= z6333_assgn63332;
        z6333_assgn63334 <= z6333_assgn63333;
        z2705_assgn2705 <= z6333_assgn63334;
        z6343_assgn63430 <= z6343_assgn6343;
        z6343_assgn63431 <= z6343_assgn63430;
        z6343_assgn63432 <= z6343_assgn63431;
        z6343_assgn63433 <= z6343_assgn63432;
        z6343_assgn63434 <= z6343_assgn63433;
        z2713_assgn2713 <= z6343_assgn63434;
        z6349_assgn63490 <= z6349_assgn6349;
        z6349_assgn63491 <= z6349_assgn63490;
        z6349_assgn63492 <= z6349_assgn63491;
        z6349_assgn63493 <= z6349_assgn63492;
        z6349_assgn63494 <= z6349_assgn63493;
        z2717_assgn2717 <= z6349_assgn63494;
        z6355_assgn63550 <= z6355_assgn6355;
        z6355_assgn63551 <= z6355_assgn63550;
        z6355_assgn63552 <= z6355_assgn63551;
        z6355_assgn63553 <= z6355_assgn63552;
        z6355_assgn63554 <= z6355_assgn63553;
        z2721_assgn2721 <= z6355_assgn63554;
        z6365_assgn63650 <= z6365_assgn6365;
        z6365_assgn63651 <= z6365_assgn63650;
        z6365_assgn63652 <= z6365_assgn63651;
        z6365_assgn63653 <= z6365_assgn63652;
        z6365_assgn63654 <= z6365_assgn63653;
        z2729_assgn2729 <= z6365_assgn63654;
        z6371_assgn63710 <= z6371_assgn6371;
        z6371_assgn63711 <= z6371_assgn63710;
        z6371_assgn63712 <= z6371_assgn63711;
        z6371_assgn63713 <= z6371_assgn63712;
        z6371_assgn63714 <= z6371_assgn63713;
        z2733_assgn2733 <= z6371_assgn63714;
        z6377_assgn63770 <= z6377_assgn6377;
        z6377_assgn63771 <= z6377_assgn63770;
        z6377_assgn63772 <= z6377_assgn63771;
        z6377_assgn63773 <= z6377_assgn63772;
        z6377_assgn63774 <= z6377_assgn63773;
        z2737_assgn2737 <= z6377_assgn63774;
        z6387_assgn63870 <= z6387_assgn6387;
        z6387_assgn63871 <= z6387_assgn63870;
        z6387_assgn63872 <= z6387_assgn63871;
        z6387_assgn63873 <= z6387_assgn63872;
        z6387_assgn63874 <= z6387_assgn63873;
        z2745_assgn2745 <= z6387_assgn63874;
        z6393_assgn63930 <= z6393_assgn6393;
        z6393_assgn63931 <= z6393_assgn63930;
        z6393_assgn63932 <= z6393_assgn63931;
        z6393_assgn63933 <= z6393_assgn63932;
        z6393_assgn63934 <= z6393_assgn63933;
        z2749_assgn2749 <= z6393_assgn63934;
        z6399_assgn63990 <= z6399_assgn6399;
        z6399_assgn63991 <= z6399_assgn63990;
        z6399_assgn63992 <= z6399_assgn63991;
        z6399_assgn63993 <= z6399_assgn63992;
        z6399_assgn63994 <= z6399_assgn63993;
        z2753_assgn2753 <= z6399_assgn63994;
        z6409_assgn64090 <= z6409_assgn6409;
        z6409_assgn64091 <= z6409_assgn64090;
        z6409_assgn64092 <= z6409_assgn64091;
        z6409_assgn64093 <= z6409_assgn64092;
        z6409_assgn64094 <= z6409_assgn64093;
        z2761_assgn2761 <= z6409_assgn64094;
        z6419_assgn64190 <= z6419_assgn6419;
        z6419_assgn64191 <= z6419_assgn64190;
        z6419_assgn64192 <= z6419_assgn64191;
        z6419_assgn64193 <= z6419_assgn64192;
        z6419_assgn64194 <= z6419_assgn64193;
        z2769_assgn2769 <= z6419_assgn64194;
        z6427_assgn64270 <= z6427_assgn6427;
        z6427_assgn64271 <= z6427_assgn64270;
        z6427_assgn64272 <= z6427_assgn64271;
        z6427_assgn64273 <= z6427_assgn64272;
        z6427_assgn64274 <= z6427_assgn64273;
        z2775_assgn2775 <= z6427_assgn64274;
        z6431_assgn64310 <= z6431_assgn6431;
        z6431_assgn64311 <= z6431_assgn64310;
        z6431_assgn64312 <= z6431_assgn64311;
        z6431_assgn64313 <= z6431_assgn64312;
        z6431_assgn64314 <= z6431_assgn64313;
        z2778_assgn2778 <= z6431_assgn64314;
        z6437_assgn64370 <= z6437_assgn6437;
        z6437_assgn64371 <= z6437_assgn64370;
        z6437_assgn64372 <= z6437_assgn64371;
        z6437_assgn64373 <= z6437_assgn64372;
        z6437_assgn64374 <= z6437_assgn64373;
        z2781_assgn2781 <= z6437_assgn64374;
        z6443_assgn64430 <= z6443_assgn6443;
        z6443_assgn64431 <= z6443_assgn64430;
        z6443_assgn64432 <= z6443_assgn64431;
        z6443_assgn64433 <= z6443_assgn64432;
        z6443_assgn64434 <= z6443_assgn64433;
        z2785_assgn2785 <= z6443_assgn64434;
        z6449_assgn64490 <= z6449_assgn6449;
        z6449_assgn64491 <= z6449_assgn64490;
        z6449_assgn64492 <= z6449_assgn64491;
        z6449_assgn64493 <= z6449_assgn64492;
        z6449_assgn64494 <= z6449_assgn64493;
        z2789_assgn2789 <= z6449_assgn64494;
        z6459_assgn64590 <= z6459_assgn6459;
        z6459_assgn64591 <= z6459_assgn64590;
        z6459_assgn64592 <= z6459_assgn64591;
        z6459_assgn64593 <= z6459_assgn64592;
        z6459_assgn64594 <= z6459_assgn64593;
        z2797_assgn2797 <= z6459_assgn64594;
        z6465_assgn64650 <= z6465_assgn6465;
        z6465_assgn64651 <= z6465_assgn64650;
        z6465_assgn64652 <= z6465_assgn64651;
        z6465_assgn64653 <= z6465_assgn64652;
        z6465_assgn64654 <= z6465_assgn64653;
        z2801_assgn2801 <= z6465_assgn64654;
        z6471_assgn64710 <= z6471_assgn6471;
        z6471_assgn64711 <= z6471_assgn64710;
        z6471_assgn64712 <= z6471_assgn64711;
        z6471_assgn64713 <= z6471_assgn64712;
        z6471_assgn64714 <= z6471_assgn64713;
        z2805_assgn2805 <= z6471_assgn64714;
        z6481_assgn64810 <= z6481_assgn6481;
        z6481_assgn64811 <= z6481_assgn64810;
        z6481_assgn64812 <= z6481_assgn64811;
        z6481_assgn64813 <= z6481_assgn64812;
        z6481_assgn64814 <= z6481_assgn64813;
        z2813_assgn2813 <= z6481_assgn64814;
        z6487_assgn64870 <= z6487_assgn6487;
        z6487_assgn64871 <= z6487_assgn64870;
        z6487_assgn64872 <= z6487_assgn64871;
        z6487_assgn64873 <= z6487_assgn64872;
        z6487_assgn64874 <= z6487_assgn64873;
        z2817_assgn2817 <= z6487_assgn64874;
        z6493_assgn64930 <= z6493_assgn6493;
        z6493_assgn64931 <= z6493_assgn64930;
        z6493_assgn64932 <= z6493_assgn64931;
        z6493_assgn64933 <= z6493_assgn64932;
        z6493_assgn64934 <= z6493_assgn64933;
        z2821_assgn2821 <= z6493_assgn64934;
        z6503_assgn65030 <= z6503_assgn6503;
        z6503_assgn65031 <= z6503_assgn65030;
        z6503_assgn65032 <= z6503_assgn65031;
        z6503_assgn65033 <= z6503_assgn65032;
        z6503_assgn65034 <= z6503_assgn65033;
        z2829_assgn2829 <= z6503_assgn65034;
        z6509_assgn65090 <= z6509_assgn6509;
        z6509_assgn65091 <= z6509_assgn65090;
        z6509_assgn65092 <= z6509_assgn65091;
        z6509_assgn65093 <= z6509_assgn65092;
        z6509_assgn65094 <= z6509_assgn65093;
        z2833_assgn2833 <= z6509_assgn65094;
        z6515_assgn65150 <= z6515_assgn6515;
        z6515_assgn65151 <= z6515_assgn65150;
        z6515_assgn65152 <= z6515_assgn65151;
        z6515_assgn65153 <= z6515_assgn65152;
        z6515_assgn65154 <= z6515_assgn65153;
        z2837_assgn2837 <= z6515_assgn65154;
        z6525_assgn65250 <= z6525_assgn6525;
        z6525_assgn65251 <= z6525_assgn65250;
        z6525_assgn65252 <= z6525_assgn65251;
        z6525_assgn65253 <= z6525_assgn65252;
        z6525_assgn65254 <= z6525_assgn65253;
        z2845_assgn2845 <= z6525_assgn65254;
        z6531_assgn65310 <= z6531_assgn6531;
        z6531_assgn65311 <= z6531_assgn65310;
        z6531_assgn65312 <= z6531_assgn65311;
        z6531_assgn65313 <= z6531_assgn65312;
        z6531_assgn65314 <= z6531_assgn65313;
        z2849_assgn2849 <= z6531_assgn65314;
        z6537_assgn65370 <= z6537_assgn6537;
        z6537_assgn65371 <= z6537_assgn65370;
        z6537_assgn65372 <= z6537_assgn65371;
        z6537_assgn65373 <= z6537_assgn65372;
        z6537_assgn65374 <= z6537_assgn65373;
        z2853_assgn2853 <= z6537_assgn65374;
        z6547_assgn65470 <= z6547_assgn6547;
        z6547_assgn65471 <= z6547_assgn65470;
        z6547_assgn65472 <= z6547_assgn65471;
        z6547_assgn65473 <= z6547_assgn65472;
        z6547_assgn65474 <= z6547_assgn65473;
        z2861_assgn2861 <= z6547_assgn65474;
        z6553_assgn65530 <= z6553_assgn6553;
        z6553_assgn65531 <= z6553_assgn65530;
        z6553_assgn65532 <= z6553_assgn65531;
        z6553_assgn65533 <= z6553_assgn65532;
        z6553_assgn65534 <= z6553_assgn65533;
        z2865_assgn2865 <= z6553_assgn65534;
        z6559_assgn65590 <= z6559_assgn6559;
        z6559_assgn65591 <= z6559_assgn65590;
        z6559_assgn65592 <= z6559_assgn65591;
        z6559_assgn65593 <= z6559_assgn65592;
        z6559_assgn65594 <= z6559_assgn65593;
        z2869_assgn2869 <= z6559_assgn65594;
        z6569_assgn65690 <= z6569_assgn6569;
        z6569_assgn65691 <= z6569_assgn65690;
        z6569_assgn65692 <= z6569_assgn65691;
        z6569_assgn65693 <= z6569_assgn65692;
        z6569_assgn65694 <= z6569_assgn65693;
        z2877_assgn2877 <= z6569_assgn65694;
        z6575_assgn65750 <= z6575_assgn6575;
        z6575_assgn65751 <= z6575_assgn65750;
        z6575_assgn65752 <= z6575_assgn65751;
        z6575_assgn65753 <= z6575_assgn65752;
        z6575_assgn65754 <= z6575_assgn65753;
        z2881_assgn2881 <= z6575_assgn65754;
        z6581_assgn65810 <= z6581_assgn6581;
        z6581_assgn65811 <= z6581_assgn65810;
        z6581_assgn65812 <= z6581_assgn65811;
        z6581_assgn65813 <= z6581_assgn65812;
        z6581_assgn65814 <= z6581_assgn65813;
        z2885_assgn2885 <= z6581_assgn65814;
        z6591_assgn65910 <= z6591_assgn6591;
        z6591_assgn65911 <= z6591_assgn65910;
        z6591_assgn65912 <= z6591_assgn65911;
        z6591_assgn65913 <= z6591_assgn65912;
        z6591_assgn65914 <= z6591_assgn65913;
        z2893_assgn2893 <= z6591_assgn65914;
        z6597_assgn65970 <= z6597_assgn6597;
        z6597_assgn65971 <= z6597_assgn65970;
        z6597_assgn65972 <= z6597_assgn65971;
        z6597_assgn65973 <= z6597_assgn65972;
        z6597_assgn65974 <= z6597_assgn65973;
        z2897_assgn2897 <= z6597_assgn65974;
        y0 <= (t6 ^ z2897_assgn2897);
        y1 <= t7;
    end

endmodule

