module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1
);
//input [31:0]S
    input clk;
    input [31:0]  t0;
    input [31:0]  t1;
    input [31:0]  r0;
    input [31:0]  r1;
    input [31:0]  r2;
    input [31:0]  r3;
    input [31:0]  r4;
    input [31:0]  r5;
    input [31:0]  dec_0;
    input [31:0]  dec_1;
    input [31:0]  dec_255;
    input [31:0]  dec_169;
    input [31:0]  dec_129;
    input [31:0]  dec_9;
    input [31:0]  dec_72;
    input [31:0]  dec_242;
    input [31:0]  dec_243;
    input [31:0]  dec_152;
    input [31:0]  dec_240;
    input [31:0]  dec_4;
    input [31:0]  dec_15;
    input [31:0]  dec_12;
    input [31:0]  dec_2;
    input [31:0]  dec_3;
    input [31:0]  dec_16;
    input [31:0]  dec_36;
    input [31:0]  dec_220;
    input [31:0]  dec_11;
    input [31:0]  dec_158;
    input [31:0]  dec_45;
    input [31:0]  dec_88;
    input [31:0]  dec_99;
//OUTPUTS
    output reg [31:0] y0;
    output reg [31:0] y1;
//Intermediate values
    wire [31:0] dec_99_inp;
    wire [31:0] dec_88_inp;
    wire [31:0] dec_45_inp;
    wire [31:0] dec_158_inp;
    wire [31:0] dec_11_inp;
    wire [31:0] dec_220_inp;
    wire [31:0] dec_36_inp;
    wire [31:0] dec_16_inp;
    wire [31:0] dec_3_inp;
    wire [31:0] dec_2_inp;
    wire [31:0] dec_12_inp;
    wire [31:0] dec_15_inp;
    wire [31:0] dec_4_inp;
    wire [31:0] dec_240_inp;
    wire [31:0] dec_152_inp;
    wire [31:0] dec_243_inp;
    wire [31:0] dec_242_inp;
    wire [31:0] dec_72_inp;
    wire [31:0] dec_9_inp;
    wire [31:0] dec_129_inp;
    wire [31:0] dec_169_inp;
    wire [31:0] dec_255_inp;
    wire [31:0] dec_1_inp;
    wire [31:0] dec_0_inp;
    wire [31:0] t0_inp;
    wire [31:0] t1_inp;
    wire [31:0] r0_inp;
    wire [31:0] r1_inp;
    wire [31:0] r2_inp;
    wire [31:0] r3_inp;
    wire [31:0] r4_inp;
    wire [31:0] r5_inp;
    wire [31:0] y_G256_newbasis0;
    wire [31:0] tempy1_G256_newbasis0;
    wire [31:0] cond1_G256_newbasis0;
    wire [31:0] negCond1_G256_newbasis0;
    wire [31:0] yxorb1_G256_newbasis0;
    wire [31:0] ny1_G256_newbasis0;
    wire [31:0] tempyIntoNegCond1_G256_newbasis0;
    wire [31:0] y1_G256_newbasis0;
    wire [31:0] x1_G256_newbasis0;
    wire [31:0] tempy2_G256_newbasis0;
    wire [31:0] cond2_G256_newbasis0;
    wire [31:0] negCond2_G256_newbasis0;
    wire [31:0] yxorb2_G256_newbasis0;
    wire [31:0] ny2_G256_newbasis0;
    wire [31:0] tempyIntoNegCond2_G256_newbasis0;
    wire [31:0] y2_G256_newbasis0;
    wire [31:0] x2_G256_newbasis0;
    wire [31:0] tempy3_G256_newbasis0;
    wire [31:0] cond3_G256_newbasis0;
    wire [31:0] negCond3_G256_newbasis0;
    wire [31:0] yxorb3_G256_newbasis0;
    wire [31:0] ny3_G256_newbasis0;
    wire [31:0] tempyIntoNegCond3_G256_newbasis0;
    wire [31:0] y3_G256_newbasis0;
    wire [31:0] x3_G256_newbasis0;
    wire [31:0] tempy4_G256_newbasis0;
    wire [31:0] cond4_G256_newbasis0;
    wire [31:0] negCond4_G256_newbasis0;
    wire [31:0] yxorb4_G256_newbasis0;
    wire [31:0] ny4_G256_newbasis0;
    wire [31:0] tempyIntoNegCond4_G256_newbasis0;
    wire [31:0] y4_G256_newbasis0;
    wire [31:0] x4_G256_newbasis0;
    wire [31:0] tempy5_G256_newbasis0;
    wire [31:0] cond5_G256_newbasis0;
    wire [31:0] negCond5_G256_newbasis0;
    wire [31:0] yxorb5_G256_newbasis0;
    wire [31:0] ny5_G256_newbasis0;
    wire [31:0] tempyIntoNegCond5_G256_newbasis0;
    wire [31:0] y5_G256_newbasis0;
    wire [31:0] x5_G256_newbasis0;
    wire [31:0] tempy6_G256_newbasis0;
    wire [31:0] cond6_G256_newbasis0;
    wire [31:0] negCond6_G256_newbasis0;
    wire [31:0] yxorb6_G256_newbasis0;
    wire [31:0] ny6_G256_newbasis0;
    wire [31:0] tempyIntoNegCond6_G256_newbasis0;
    wire [31:0] y6_G256_newbasis0;
    wire [31:0] x6_G256_newbasis0;
    wire [31:0] tempy7_G256_newbasis0;
    wire [31:0] cond7_G256_newbasis0;
    wire [31:0] negCond7_G256_newbasis0;
    wire [31:0] yxorb7_G256_newbasis0;
    wire [31:0] ny7_G256_newbasis0;
    wire [31:0] tempyIntoNegCond7_G256_newbasis0;
    wire [31:0] y7_G256_newbasis0;
    wire [31:0] x7_G256_newbasis0;
    wire [31:0] tempy8_G256_newbasis0;
    wire [31:0] cond8_G256_newbasis0;
    wire [31:0] negCond8_G256_newbasis0;
    wire [31:0] yxorb8_G256_newbasis0;
    wire [31:0] ny8_G256_newbasis0;
    wire [31:0] tempyIntoNegCond8_G256_newbasis0;
    wire [31:0] y8_G256_newbasis0;
    wire [31:0] z3873_assgn3873;
    reg [31:0] z3873_assgn38730;
    reg [31:0] z3873_assgn38731;
    reg [31:0] z3873_assgn38732;
    reg [31:0] z3873_assgn38733;
    reg [31:0] z3873_assgn38734;
    reg [31:0] z3873_assgn38735;
    reg [31:0] z3873_assgn38736;
    reg [31:0] z3873_assgn38737;
    reg [31:0] z3873_assgn38738;
    reg [31:0] z3873_assgn38739;
    reg [31:0] z3873_assgn387310;
    reg [31:0] x8_G256_newbasis0;
    wire [31:0] t2;
    wire [31:0] z_y_G256_newbasis0;
    wire [31:0] z_tempy1_G256_newbasis0;
    wire [31:0] z_cond1_G256_newbasis0;
    wire [31:0] z_negCond1_G256_newbasis0;
    wire [31:0] z_yxorb1_G256_newbasis0;
    wire [31:0] z_ny1_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond1_G256_newbasis0;
    wire [31:0] z_y1_G256_newbasis0;
    wire [31:0] z_x1_G256_newbasis0;
    wire [31:0] z_tempy2_G256_newbasis0;
    wire [31:0] z_cond2_G256_newbasis0;
    wire [31:0] z_negCond2_G256_newbasis0;
    wire [31:0] z_yxorb2_G256_newbasis0;
    wire [31:0] z_ny2_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond2_G256_newbasis0;
    wire [31:0] z_y2_G256_newbasis0;
    wire [31:0] z_x2_G256_newbasis0;
    wire [31:0] z_tempy3_G256_newbasis0;
    wire [31:0] z_cond3_G256_newbasis0;
    wire [31:0] z_negCond3_G256_newbasis0;
    wire [31:0] z_yxorb3_G256_newbasis0;
    wire [31:0] z_ny3_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond3_G256_newbasis0;
    wire [31:0] z_y3_G256_newbasis0;
    wire [31:0] z_x3_G256_newbasis0;
    wire [31:0] z_tempy4_G256_newbasis0;
    wire [31:0] z_cond4_G256_newbasis0;
    wire [31:0] z_negCond4_G256_newbasis0;
    wire [31:0] z_yxorb4_G256_newbasis0;
    wire [31:0] z_ny4_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond4_G256_newbasis0;
    wire [31:0] z_y4_G256_newbasis0;
    wire [31:0] z_x4_G256_newbasis0;
    wire [31:0] z_tempy5_G256_newbasis0;
    wire [31:0] z_cond5_G256_newbasis0;
    wire [31:0] z_negCond5_G256_newbasis0;
    wire [31:0] z_yxorb5_G256_newbasis0;
    wire [31:0] z_ny5_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond5_G256_newbasis0;
    wire [31:0] z_y5_G256_newbasis0;
    wire [31:0] z_x5_G256_newbasis0;
    wire [31:0] z_tempy6_G256_newbasis0;
    wire [31:0] z_cond6_G256_newbasis0;
    wire [31:0] z_negCond6_G256_newbasis0;
    wire [31:0] z_yxorb6_G256_newbasis0;
    wire [31:0] z_ny6_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond6_G256_newbasis0;
    wire [31:0] z_y6_G256_newbasis0;
    wire [31:0] z_x6_G256_newbasis0;
    wire [31:0] z_tempy7_G256_newbasis0;
    wire [31:0] z_cond7_G256_newbasis0;
    wire [31:0] z_negCond7_G256_newbasis0;
    wire [31:0] z_yxorb7_G256_newbasis0;
    wire [31:0] z_ny7_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond7_G256_newbasis0;
    wire [31:0] z_y7_G256_newbasis0;
    wire [31:0] z_x7_G256_newbasis0;
    wire [31:0] z_tempy8_G256_newbasis0;
    wire [31:0] z_cond8_G256_newbasis0;
    wire [31:0] z_negCond8_G256_newbasis0;
    wire [31:0] z_yxorb8_G256_newbasis0;
    wire [31:0] z_ny8_G256_newbasis0;
    wire [31:0] z_tempyIntoNegCond8_G256_newbasis0;
    wire [31:0] z_y8_G256_newbasis0;
    wire [31:0] z4005_assgn4005;
    reg [31:0] z4005_assgn40050;
    reg [31:0] z4005_assgn40051;
    reg [31:0] z4005_assgn40052;
    reg [31:0] z4005_assgn40053;
    reg [31:0] z4005_assgn40054;
    reg [31:0] z4005_assgn40055;
    reg [31:0] z4005_assgn40056;
    reg [31:0] z4005_assgn40057;
    reg [31:0] z4005_assgn40058;
    reg [31:0] z4005_assgn40059;
    reg [31:0] z4005_assgn400510;
    reg [31:0] z_x8_G256_newbasis0;
    wire [31:0] t3;
    wire [31:0] a0_0_G256_inv0;
    wire [31:0] a1_0_G256_inv0;
    wire [31:0] a0_G256_inv0;
    wire [31:0] a1_G256_inv0;
    wire [31:0] b0_G256_inv0;
    wire [31:0] b1_G256_inv0;
    wire [31:0] a0xorb0_G256_inv0;
    wire [31:0] a1xorb1_G256_inv0;
    wire [31:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_G16_sq_scl0_G256_inv0;
    wire [31:0] b0_G16_sq_scl0_G256_inv0;
    wire [31:0] b1_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_0_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [31:0] q0_G16_sq_scl0_G256_inv0;
    wire [31:0] q1_G16_sq_scl0_G256_inv0;
    wire [31:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [31:0] p1ls2_G16_sq_scl0_G256_inv0;
    wire [31:0] c0_G256_inv0;
    wire [31:0] c1_G256_inv0;
    wire [31:0] r00_G16_mul0_G256_inv0;
    wire [31:0] r10_G16_mul0_G256_inv0;
    wire [31:0] r20_G16_mul0_G256_inv0;
    wire [31:0] r30_G16_mul0_G256_inv0;
    wire [31:0] r40_G16_mul0_G256_inv0;
    wire [31:0] r50_G16_mul0_G256_inv0;
    wire [31:0] a0_0_G16_mul0_G256_inv0;
    wire [31:0] a1_0_G16_mul0_G256_inv0;
    wire [31:0] a0_G16_mul0_G256_inv0;
    wire [31:0] a1_G16_mul0_G256_inv0;
    wire [31:0] b0_G16_mul0_G256_inv0;
    wire [31:0] b1_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G16_mul0_G256_inv0;
    wire [31:0] c0_G16_mul0_G256_inv0;
    wire [31:0] c1_G16_mul0_G256_inv0;
    wire [31:0] d0_G16_mul0_G256_inv0;
    wire [31:0] d1_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G16_mul0_G256_inv0;
    wire [31:0] cxord_0_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G16_mul0_G256_inv0;
    wire [31:0] cxord_1_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r30_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r40_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r50_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] a1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] b1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] cxord_1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m3_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m3_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p4_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i1_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i0_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar0_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] e0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] e1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m3_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m3_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p4_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i1_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i0_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar1_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] m3_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] m3_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p4_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i1_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] i0_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar2_G4_mul0_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0;
    reg [31:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] z4371_assgn4371;
    reg [31:0] z4371_assgn43710;
    reg [31:0] z4371_assgn43711;
    reg [31:0] z691_assgn691;
    wire [31:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [31:0] e0_G16_mul0_G256_inv0;
    wire [31:0] e1_G16_mul0_G256_inv0;
    wire [31:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z4381_assgn4381;
    reg [31:0] z4381_assgn43810;
    reg [31:0] z4381_assgn43811;
    reg [31:0] z699_assgn699;
    wire [31:0] a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z4387_assgn4387;
    reg [31:0] z4387_assgn43870;
    reg [31:0] z4387_assgn43871;
    reg [31:0] z703_assgn703;
    wire [31:0] a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z4393_assgn4393;
    reg [31:0] z4393_assgn43930;
    reg [31:0] z4393_assgn43931;
    reg [31:0] z707_assgn707;
    wire [31:0] b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] z4405_assgn4405;
    reg [31:0] z4405_assgn44050;
    reg [31:0] z4405_assgn44051;
    reg [31:0] z717_assgn717;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [31:0] e01_G16_mul0_G256_inv0;
    wire [31:0] e11_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r30_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r40_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r50_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] a1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] b1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m3_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m3_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p4_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i1_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i0_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar0_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] e0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] e1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m3_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m3_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p4_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i1_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i0_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar1_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] m3_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] m3_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p4_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i1_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] i0_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar2_G4_mul1_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0;
    reg [31:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] z4625_assgn4625;
    reg [31:0] z4625_assgn46250;
    reg [31:0] z4625_assgn46251;
    reg [31:0] z935_assgn935;
    wire [31:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [31:0] p0_0_G16_mul0_G256_inv0;
    wire [31:0] p1_0_G16_mul0_G256_inv0;
    wire [31:0] p0_G16_mul0_G256_inv0;
    wire [31:0] p1_G16_mul0_G256_inv0;
    wire [31:0] r00_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r10_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r20_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r30_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r40_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r50_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] a1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] b1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] c1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] d1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m3_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m3_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p4_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i1_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i0_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar0_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] e0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] e1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m3_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m3_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p4_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i1_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i0_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar1_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] m3_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] m3_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p4_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r2_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i2_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] r3_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i3_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i1_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i2_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] i0_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    reg [31:0] i3_comar2_G4_mul2_G16_mul0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0;
    reg [31:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] z4847_assgn4847;
    reg [31:0] z4847_assgn48470;
    reg [31:0] z4847_assgn48471;
    reg [31:0] z1155_assgn1155;
    wire [31:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [31:0] q0_0_G16_mul0_G256_inv0;
    wire [31:0] q1_0_G16_mul0_G256_inv0;
    wire [31:0] q0_G16_mul0_G256_inv0;
    wire [31:0] q1_G16_mul0_G256_inv0;
    wire [31:0] p0ls2_G16_mul0_G256_inv0;
    wire [31:0] z4861_assgn4861;
    reg [31:0] z4861_assgn48610;
    reg [31:0] z4861_assgn48611;
    reg [31:0] z1167_assgn1167;
    wire [31:0] p1ls2_G16_mul0_G256_inv0;
    wire [31:0] d0_G256_inv0;
    wire [31:0] d1_G256_inv0;
    wire [31:0] c0xord0_G256_inv0;
    wire [31:0] z4871_assgn4871;
    reg [31:0] z4871_assgn48710;
    reg [31:0] z4871_assgn48711;
    reg [31:0] z1176_assgn1176;
    wire [31:0] c1xord1_G256_inv0;
    wire [31:0] r00_G16_inv0_G256_inv0;
    wire [31:0] r10_G16_inv0_G256_inv0;
    wire [31:0] r20_G16_inv0_G256_inv0;
    wire [31:0] r30_G16_inv0_G256_inv0;
    wire [31:0] r40_G16_inv0_G256_inv0;
    wire [31:0] r50_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G16_inv0_G256_inv0;
    wire [31:0] z4889_assgn4889;
    reg [31:0] z4889_assgn48890;
    reg [31:0] z4889_assgn48891;
    reg [31:0] z1191_assgn1191;
    wire [31:0] a1_0_G16_inv0_G256_inv0;
    wire [31:0] a0_G16_inv0_G256_inv0;
    wire [31:0] z4895_assgn4895;
    reg [31:0] z4895_assgn48950;
    reg [31:0] z4895_assgn48951;
    reg [31:0] z1195_assgn1195;
    wire [31:0] a1_G16_inv0_G256_inv0;
    wire [31:0] b0_G16_inv0_G256_inv0;
    wire [31:0] z4901_assgn4901;
    reg [31:0] z4901_assgn49010;
    reg [31:0] z4901_assgn49011;
    reg [31:0] z1199_assgn1199;
    wire [31:0] b1_G16_inv0_G256_inv0;
    wire [31:0] a0xorb0_G16_inv0_G256_inv0;
    wire [31:0] a1xorb1_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4911_assgn4911;
    reg [31:0] z4911_assgn49110;
    reg [31:0] z4911_assgn49111;
    reg [31:0] z1207_assgn1207;
    wire [31:0] a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4917_assgn4917;
    reg [31:0] z4917_assgn49170;
    reg [31:0] z4917_assgn49171;
    reg [31:0] z1211_assgn1211;
    wire [31:0] a1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4923_assgn4923;
    reg [31:0] z4923_assgn49230;
    reg [31:0] z4923_assgn49231;
    reg [31:0] z1215_assgn1215;
    wire [31:0] b1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] z4929_assgn4929;
    reg [31:0] z4929_assgn49290;
    reg [31:0] z4929_assgn49291;
    reg [31:0] z1219_assgn1219;
    wire [31:0] b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [31:0] c0_0_G16_inv0_G256_inv0;
    wire [31:0] c1_0_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4939_assgn4939;
    reg [31:0] z4939_assgn49390;
    reg [31:0] z4939_assgn49391;
    reg [31:0] z1227_assgn1227;
    wire [31:0] a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4945_assgn4945;
    reg [31:0] z4945_assgn49450;
    reg [31:0] z4945_assgn49451;
    reg [31:0] z1231_assgn1231;
    wire [31:0] a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4951_assgn4951;
    reg [31:0] z4951_assgn49510;
    reg [31:0] z4951_assgn49511;
    reg [31:0] z1235_assgn1235;
    wire [31:0] b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] z4963_assgn4963;
    reg [31:0] z4963_assgn49630;
    reg [31:0] z4963_assgn49631;
    reg [31:0] z1245_assgn1245;
    wire [31:0] p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [31:0] c0_G16_inv0_G256_inv0;
    wire [31:0] c1_G16_inv0_G256_inv0;
    wire [31:0] r00_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r10_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r20_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r30_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r40_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r50_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4987_assgn4987;
    reg [31:0] z4987_assgn49870;
    reg [31:0] z4987_assgn49871;
    reg [31:0] z1267_assgn1267;
    wire [31:0] a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4993_assgn4993;
    reg [31:0] z4993_assgn49930;
    reg [31:0] z4993_assgn49931;
    reg [31:0] z1271_assgn1271;
    wire [31:0] a1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z4999_assgn4999;
    reg [31:0] z4999_assgn49990;
    reg [31:0] z4999_assgn49991;
    reg [31:0] z1275_assgn1275;
    wire [31:0] b1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5005_assgn5005;
    reg [31:0] z5005_assgn50050;
    reg [31:0] z5005_assgn50051;
    reg [31:0] z1279_assgn1279;
    wire [31:0] c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5011_assgn5011;
    reg [31:0] z5011_assgn50110;
    reg [31:0] z5011_assgn50111;
    reg [31:0] z1283_assgn1283;
    wire [31:0] c1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5017_assgn5017;
    reg [31:0] z5017_assgn50170;
    reg [31:0] z5017_assgn50171;
    reg [31:0] z1287_assgn1287;
    wire [31:0] d1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5043_assgn5043;
    reg [31:0] z5043_assgn50430;
    reg [31:0] z5043_assgn50431;
    reg [31:0] z1311_assgn1311;
    wire [31:0] m1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5049_assgn5049;
    reg [31:0] z5049_assgn50490;
    reg [31:0] z5049_assgn50491;
    reg [31:0] z1315_assgn1315;
    wire [31:0] m3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5053_assgn5053;
    reg [31:0] z5053_assgn50530;
    reg [31:0] z5053_assgn50531;
    reg [31:0] z5053_assgn50532;
    reg [31:0] z1318_assgn1318;
    reg [31:0] m1_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5057_assgn5057;
    reg [31:0] z5057_assgn50570;
    reg [31:0] z5057_assgn50571;
    reg [31:0] z5057_assgn50572;
    reg [31:0] z1319_assgn1319;
    reg [31:0] m3_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p4_comar0_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5067_assgn5067;
    reg [31:0] z5067_assgn50670;
    reg [31:0] z5067_assgn50671;
    reg [31:0] z5067_assgn50672;
    reg [31:0] z1327_assgn1327;
    wire [31:0] i1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5071_assgn5071;
    reg [31:0] z5071_assgn50710;
    reg [31:0] z5071_assgn50711;
    reg [31:0] z5071_assgn50712;
    reg [31:0] z1329_assgn1329;
    wire [31:0] i2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5075_assgn5075;
    reg [31:0] z5075_assgn50750;
    reg [31:0] z5075_assgn50751;
    reg [31:0] z5075_assgn50752;
    reg [31:0] z1331_assgn1331;
    wire [31:0] i3_comar0_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] i1_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] i2_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5081_assgn5081;
    reg [31:0] z5081_assgn50810;
    reg [31:0] z5081_assgn50811;
    reg [31:0] z5081_assgn50812;
    reg [31:0] z1336_assgn1336;
    reg [31:0] i3_comar0_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] e0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] e1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5111_assgn5111;
    reg [31:0] z5111_assgn51110;
    reg [31:0] z5111_assgn51111;
    reg [31:0] z1363_assgn1363;
    wire [31:0] m1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5117_assgn5117;
    reg [31:0] z5117_assgn51170;
    reg [31:0] z5117_assgn51171;
    reg [31:0] z1367_assgn1367;
    wire [31:0] m3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5121_assgn5121;
    reg [31:0] z5121_assgn51210;
    reg [31:0] z5121_assgn51211;
    reg [31:0] z5121_assgn51212;
    reg [31:0] z1370_assgn1370;
    reg [31:0] m1_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5125_assgn5125;
    reg [31:0] z5125_assgn51250;
    reg [31:0] z5125_assgn51251;
    reg [31:0] z5125_assgn51252;
    reg [31:0] z1371_assgn1371;
    reg [31:0] m3_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p4_comar1_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5135_assgn5135;
    reg [31:0] z5135_assgn51350;
    reg [31:0] z5135_assgn51351;
    reg [31:0] z5135_assgn51352;
    reg [31:0] z1379_assgn1379;
    wire [31:0] i1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5139_assgn5139;
    reg [31:0] z5139_assgn51390;
    reg [31:0] z5139_assgn51391;
    reg [31:0] z5139_assgn51392;
    reg [31:0] z1381_assgn1381;
    wire [31:0] i2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5143_assgn5143;
    reg [31:0] z5143_assgn51430;
    reg [31:0] z5143_assgn51431;
    reg [31:0] z5143_assgn51432;
    reg [31:0] z1383_assgn1383;
    wire [31:0] i3_comar1_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] i1_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] i2_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5149_assgn5149;
    reg [31:0] z5149_assgn51490;
    reg [31:0] z5149_assgn51491;
    reg [31:0] z5149_assgn51492;
    reg [31:0] z1388_assgn1388;
    reg [31:0] i3_comar1_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5183_assgn5183;
    reg [31:0] z5183_assgn51830;
    reg [31:0] z5183_assgn51831;
    reg [31:0] z1419_assgn1419;
    wire [31:0] m1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5189_assgn5189;
    reg [31:0] z5189_assgn51890;
    reg [31:0] z5189_assgn51891;
    reg [31:0] z1423_assgn1423;
    wire [31:0] m3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5193_assgn5193;
    reg [31:0] z5193_assgn51930;
    reg [31:0] z5193_assgn51931;
    reg [31:0] z5193_assgn51932;
    reg [31:0] z1426_assgn1426;
    reg [31:0] m1_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5197_assgn5197;
    reg [31:0] z5197_assgn51970;
    reg [31:0] z5197_assgn51971;
    reg [31:0] z5197_assgn51972;
    reg [31:0] z1427_assgn1427;
    reg [31:0] m3_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p4_comar2_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5207_assgn5207;
    reg [31:0] z5207_assgn52070;
    reg [31:0] z5207_assgn52071;
    reg [31:0] z5207_assgn52072;
    reg [31:0] z1435_assgn1435;
    wire [31:0] i1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5211_assgn5211;
    reg [31:0] z5211_assgn52110;
    reg [31:0] z5211_assgn52111;
    reg [31:0] z5211_assgn52112;
    reg [31:0] z1437_assgn1437;
    wire [31:0] i2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5215_assgn5215;
    reg [31:0] z5215_assgn52150;
    reg [31:0] z5215_assgn52151;
    reg [31:0] z5215_assgn52152;
    reg [31:0] z1439_assgn1439;
    wire [31:0] i3_comar2_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] i1_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    reg [31:0] i2_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5221_assgn5221;
    reg [31:0] z5221_assgn52210;
    reg [31:0] z5221_assgn52211;
    reg [31:0] z5221_assgn52212;
    reg [31:0] z1444_assgn1444;
    reg [31:0] i3_comar2_G4_mul3_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0;
    reg [31:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] z5243_assgn5243;
    reg [31:0] z5243_assgn52430;
    reg [31:0] z5243_assgn52431;
    reg [31:0] z5243_assgn52432;
    reg [31:0] z5243_assgn52433;
    reg [31:0] z5243_assgn52434;
    reg [31:0] z1463_assgn1463;
    wire [31:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [31:0] d0_G16_inv0_G256_inv0;
    wire [31:0] d1_G16_inv0_G256_inv0;
    wire [31:0] c0xord0_G16_inv0_G256_inv0;
    wire [31:0] z5253_assgn5253;
    reg [31:0] z5253_assgn52530;
    reg [31:0] z5253_assgn52531;
    reg [31:0] z1472_assgn1472;
    wire [31:0] c1xord1_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z5259_assgn5259;
    reg [31:0] z5259_assgn52590;
    reg [31:0] z5259_assgn52591;
    reg [31:0] z5259_assgn52592;
    reg [31:0] z5259_assgn52593;
    reg [31:0] z5259_assgn52594;
    reg [31:0] z1475_assgn1475;
    wire [31:0] a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z5265_assgn5265;
    reg [31:0] z5265_assgn52650;
    reg [31:0] z5265_assgn52651;
    reg [31:0] z5265_assgn52652;
    reg [31:0] z5265_assgn52653;
    reg [31:0] z5265_assgn52654;
    reg [31:0] z1479_assgn1479;
    wire [31:0] a1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z5271_assgn5271;
    reg [31:0] z5271_assgn52710;
    reg [31:0] z5271_assgn52711;
    reg [31:0] z5271_assgn52712;
    reg [31:0] z5271_assgn52713;
    reg [31:0] z5271_assgn52714;
    reg [31:0] z1483_assgn1483;
    wire [31:0] b1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] z5277_assgn5277;
    reg [31:0] z5277_assgn52770;
    reg [31:0] z5277_assgn52771;
    reg [31:0] z5277_assgn52772;
    reg [31:0] z5277_assgn52773;
    reg [31:0] z5277_assgn52774;
    reg [31:0] z1487_assgn1487;
    wire [31:0] b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [31:0] e0_G16_inv0_G256_inv0;
    wire [31:0] e1_G16_inv0_G256_inv0;
    wire [31:0] r00_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r10_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r20_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r30_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r40_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r50_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5299_assgn5299;
    reg [31:0] z5299_assgn52990;
    reg [31:0] z5299_assgn52991;
    reg [31:0] z5299_assgn52992;
    reg [31:0] z5299_assgn52993;
    reg [31:0] z5299_assgn52994;
    reg [31:0] z1507_assgn1507;
    wire [31:0] a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5305_assgn5305;
    reg [31:0] z5305_assgn53050;
    reg [31:0] z5305_assgn53051;
    reg [31:0] z5305_assgn53052;
    reg [31:0] z5305_assgn53053;
    reg [31:0] z5305_assgn53054;
    reg [31:0] z1511_assgn1511;
    wire [31:0] a1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5311_assgn5311;
    reg [31:0] z5311_assgn53110;
    reg [31:0] z5311_assgn53111;
    reg [31:0] z5311_assgn53112;
    reg [31:0] z5311_assgn53113;
    reg [31:0] z5311_assgn53114;
    reg [31:0] z1515_assgn1515;
    wire [31:0] b1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5317_assgn5317;
    reg [31:0] z5317_assgn53170;
    reg [31:0] z5317_assgn53171;
    reg [31:0] z1519_assgn1519;
    wire [31:0] c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5323_assgn5323;
    reg [31:0] z5323_assgn53230;
    reg [31:0] z5323_assgn53231;
    reg [31:0] z1523_assgn1523;
    wire [31:0] c1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5329_assgn5329;
    reg [31:0] z5329_assgn53290;
    reg [31:0] z5329_assgn53291;
    reg [31:0] z1527_assgn1527;
    wire [31:0] d1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5355_assgn5355;
    reg [31:0] z5355_assgn53550;
    reg [31:0] z5355_assgn53551;
    reg [31:0] z1551_assgn1551;
    wire [31:0] m1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5361_assgn5361;
    reg [31:0] z5361_assgn53610;
    reg [31:0] z5361_assgn53611;
    reg [31:0] z5361_assgn53612;
    reg [31:0] z5361_assgn53613;
    reg [31:0] z5361_assgn53614;
    reg [31:0] z1555_assgn1555;
    wire [31:0] m3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5365_assgn5365;
    reg [31:0] z5365_assgn53650;
    reg [31:0] z5365_assgn53651;
    reg [31:0] z5365_assgn53652;
    reg [31:0] z1558_assgn1558;
    reg [31:0] m1_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5369_assgn5369;
    reg [31:0] z5369_assgn53690;
    reg [31:0] z5369_assgn53691;
    reg [31:0] z5369_assgn53692;
    reg [31:0] z5369_assgn53693;
    reg [31:0] z5369_assgn53694;
    reg [31:0] z5369_assgn53695;
    reg [31:0] z1559_assgn1559;
    reg [31:0] m3_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5375_assgn5375;
    reg [31:0] z5375_assgn53750;
    reg [31:0] z5375_assgn53751;
    reg [31:0] z5375_assgn53752;
    reg [31:0] z1563_assgn1563;
    wire [31:0] p4_comar0_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5381_assgn5381;
    reg [31:0] z5381_assgn53810;
    reg [31:0] z5381_assgn53811;
    reg [31:0] z5381_assgn53812;
    reg [31:0] z1567_assgn1567;
    wire [31:0] i1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5385_assgn5385;
    reg [31:0] z5385_assgn53850;
    reg [31:0] z5385_assgn53851;
    reg [31:0] z5385_assgn53852;
    reg [31:0] z5385_assgn53853;
    reg [31:0] z5385_assgn53854;
    reg [31:0] z5385_assgn53855;
    reg [31:0] z1569_assgn1569;
    wire [31:0] i2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5389_assgn5389;
    reg [31:0] z5389_assgn53890;
    reg [31:0] z5389_assgn53891;
    reg [31:0] z5389_assgn53892;
    reg [31:0] z5389_assgn53893;
    reg [31:0] z5389_assgn53894;
    reg [31:0] z5389_assgn53895;
    reg [31:0] z1571_assgn1571;
    wire [31:0] i3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5393_assgn5393;
    reg [31:0] z5393_assgn53930;
    reg [31:0] z5393_assgn53931;
    reg [31:0] z5393_assgn53932;
    reg [31:0] z1574_assgn1574;
    reg [31:0] i2_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5397_assgn5397;
    reg [31:0] z5397_assgn53970;
    reg [31:0] z5397_assgn53971;
    reg [31:0] z5397_assgn53972;
    reg [31:0] z5397_assgn53973;
    reg [31:0] z5397_assgn53974;
    reg [31:0] z5397_assgn53975;
    reg [31:0] z1576_assgn1576;
    reg [31:0] i3_comar0_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] e0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] e1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5427_assgn5427;
    reg [31:0] z5427_assgn54270;
    reg [31:0] z5427_assgn54271;
    reg [31:0] z1603_assgn1603;
    wire [31:0] m1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5433_assgn5433;
    reg [31:0] z5433_assgn54330;
    reg [31:0] z5433_assgn54331;
    reg [31:0] z5433_assgn54332;
    reg [31:0] z5433_assgn54333;
    reg [31:0] z5433_assgn54334;
    reg [31:0] z1607_assgn1607;
    wire [31:0] m3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5437_assgn5437;
    reg [31:0] z5437_assgn54370;
    reg [31:0] z5437_assgn54371;
    reg [31:0] z5437_assgn54372;
    reg [31:0] z1610_assgn1610;
    reg [31:0] m1_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5441_assgn5441;
    reg [31:0] z5441_assgn54410;
    reg [31:0] z5441_assgn54411;
    reg [31:0] z5441_assgn54412;
    reg [31:0] z5441_assgn54413;
    reg [31:0] z5441_assgn54414;
    reg [31:0] z5441_assgn54415;
    reg [31:0] z1611_assgn1611;
    reg [31:0] m3_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5447_assgn5447;
    reg [31:0] z5447_assgn54470;
    reg [31:0] z5447_assgn54471;
    reg [31:0] z5447_assgn54472;
    reg [31:0] z1615_assgn1615;
    wire [31:0] p4_comar1_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5453_assgn5453;
    reg [31:0] z5453_assgn54530;
    reg [31:0] z5453_assgn54531;
    reg [31:0] z5453_assgn54532;
    reg [31:0] z1619_assgn1619;
    wire [31:0] i1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5457_assgn5457;
    reg [31:0] z5457_assgn54570;
    reg [31:0] z5457_assgn54571;
    reg [31:0] z5457_assgn54572;
    reg [31:0] z5457_assgn54573;
    reg [31:0] z5457_assgn54574;
    reg [31:0] z5457_assgn54575;
    reg [31:0] z1621_assgn1621;
    wire [31:0] i2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5461_assgn5461;
    reg [31:0] z5461_assgn54610;
    reg [31:0] z5461_assgn54611;
    reg [31:0] z5461_assgn54612;
    reg [31:0] z5461_assgn54613;
    reg [31:0] z5461_assgn54614;
    reg [31:0] z5461_assgn54615;
    reg [31:0] z1623_assgn1623;
    wire [31:0] i3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5465_assgn5465;
    reg [31:0] z5465_assgn54650;
    reg [31:0] z5465_assgn54651;
    reg [31:0] z5465_assgn54652;
    reg [31:0] z1626_assgn1626;
    reg [31:0] i2_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5469_assgn5469;
    reg [31:0] z5469_assgn54690;
    reg [31:0] z5469_assgn54691;
    reg [31:0] z5469_assgn54692;
    reg [31:0] z5469_assgn54693;
    reg [31:0] z5469_assgn54694;
    reg [31:0] z5469_assgn54695;
    reg [31:0] z1628_assgn1628;
    reg [31:0] i3_comar1_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5503_assgn5503;
    reg [31:0] z5503_assgn55030;
    reg [31:0] z5503_assgn55031;
    reg [31:0] z1659_assgn1659;
    wire [31:0] m1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5509_assgn5509;
    reg [31:0] z5509_assgn55090;
    reg [31:0] z5509_assgn55091;
    reg [31:0] z5509_assgn55092;
    reg [31:0] z5509_assgn55093;
    reg [31:0] z5509_assgn55094;
    reg [31:0] z1663_assgn1663;
    wire [31:0] m3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5513_assgn5513;
    reg [31:0] z5513_assgn55130;
    reg [31:0] z5513_assgn55131;
    reg [31:0] z5513_assgn55132;
    reg [31:0] z1666_assgn1666;
    reg [31:0] m1_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5517_assgn5517;
    reg [31:0] z5517_assgn55170;
    reg [31:0] z5517_assgn55171;
    reg [31:0] z5517_assgn55172;
    reg [31:0] z5517_assgn55173;
    reg [31:0] z5517_assgn55174;
    reg [31:0] z5517_assgn55175;
    reg [31:0] z1667_assgn1667;
    reg [31:0] m3_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5523_assgn5523;
    reg [31:0] z5523_assgn55230;
    reg [31:0] z5523_assgn55231;
    reg [31:0] z5523_assgn55232;
    reg [31:0] z1671_assgn1671;
    wire [31:0] p4_comar2_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5529_assgn5529;
    reg [31:0] z5529_assgn55290;
    reg [31:0] z5529_assgn55291;
    reg [31:0] z5529_assgn55292;
    reg [31:0] z1675_assgn1675;
    wire [31:0] i1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5533_assgn5533;
    reg [31:0] z5533_assgn55330;
    reg [31:0] z5533_assgn55331;
    reg [31:0] z5533_assgn55332;
    reg [31:0] z5533_assgn55333;
    reg [31:0] z5533_assgn55334;
    reg [31:0] z5533_assgn55335;
    reg [31:0] z1677_assgn1677;
    wire [31:0] i2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5537_assgn5537;
    reg [31:0] z5537_assgn55370;
    reg [31:0] z5537_assgn55371;
    reg [31:0] z5537_assgn55372;
    reg [31:0] z5537_assgn55373;
    reg [31:0] z5537_assgn55374;
    reg [31:0] z5537_assgn55375;
    reg [31:0] z1679_assgn1679;
    wire [31:0] i3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5541_assgn5541;
    reg [31:0] z5541_assgn55410;
    reg [31:0] z5541_assgn55411;
    reg [31:0] z5541_assgn55412;
    reg [31:0] z1682_assgn1682;
    reg [31:0] i2_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5545_assgn5545;
    reg [31:0] z5545_assgn55450;
    reg [31:0] z5545_assgn55451;
    reg [31:0] z5545_assgn55452;
    reg [31:0] z5545_assgn55453;
    reg [31:0] z5545_assgn55454;
    reg [31:0] z5545_assgn55455;
    reg [31:0] z1684_assgn1684;
    reg [31:0] i3_comar2_G4_mul4_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0;
    reg [31:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] z5567_assgn5567;
    reg [31:0] z5567_assgn55670;
    reg [31:0] z5567_assgn55671;
    reg [31:0] z5567_assgn55672;
    reg [31:0] z5567_assgn55673;
    reg [31:0] z5567_assgn55674;
    reg [31:0] z5567_assgn55675;
    reg [31:0] z5567_assgn55676;
    reg [31:0] z5567_assgn55677;
    reg [31:0] z1703_assgn1703;
    wire [31:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [31:0] p0_G16_inv0_G256_inv0;
    wire [31:0] p1_G16_inv0_G256_inv0;
    wire [31:0] r00_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r10_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r20_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r30_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r40_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r50_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5589_assgn5589;
    reg [31:0] z5589_assgn55890;
    reg [31:0] z5589_assgn55891;
    reg [31:0] z5589_assgn55892;
    reg [31:0] z5589_assgn55893;
    reg [31:0] z5589_assgn55894;
    reg [31:0] z1723_assgn1723;
    wire [31:0] a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5595_assgn5595;
    reg [31:0] z5595_assgn55950;
    reg [31:0] z5595_assgn55951;
    reg [31:0] z5595_assgn55952;
    reg [31:0] z5595_assgn55953;
    reg [31:0] z5595_assgn55954;
    reg [31:0] z1727_assgn1727;
    wire [31:0] a1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5601_assgn5601;
    reg [31:0] z5601_assgn56010;
    reg [31:0] z5601_assgn56011;
    reg [31:0] z5601_assgn56012;
    reg [31:0] z5601_assgn56013;
    reg [31:0] z5601_assgn56014;
    reg [31:0] z1731_assgn1731;
    wire [31:0] b1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5607_assgn5607;
    reg [31:0] z5607_assgn56070;
    reg [31:0] z5607_assgn56071;
    reg [31:0] z1735_assgn1735;
    wire [31:0] c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5613_assgn5613;
    reg [31:0] z5613_assgn56130;
    reg [31:0] z5613_assgn56131;
    reg [31:0] z1739_assgn1739;
    wire [31:0] c1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5619_assgn5619;
    reg [31:0] z5619_assgn56190;
    reg [31:0] z5619_assgn56191;
    reg [31:0] z1743_assgn1743;
    wire [31:0] d1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] axorb_1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r00_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m0_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5645_assgn5645;
    reg [31:0] z5645_assgn56450;
    reg [31:0] z5645_assgn56451;
    reg [31:0] z1767_assgn1767;
    wire [31:0] m1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5651_assgn5651;
    reg [31:0] z5651_assgn56510;
    reg [31:0] z5651_assgn56511;
    reg [31:0] z5651_assgn56512;
    reg [31:0] z5651_assgn56513;
    reg [31:0] z5651_assgn56514;
    reg [31:0] z1771_assgn1771;
    wire [31:0] m3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5655_assgn5655;
    reg [31:0] z5655_assgn56550;
    reg [31:0] z5655_assgn56551;
    reg [31:0] z5655_assgn56552;
    reg [31:0] z1774_assgn1774;
    reg [31:0] m1_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5659_assgn5659;
    reg [31:0] z5659_assgn56590;
    reg [31:0] z5659_assgn56591;
    reg [31:0] z5659_assgn56592;
    reg [31:0] z5659_assgn56593;
    reg [31:0] z5659_assgn56594;
    reg [31:0] z5659_assgn56595;
    reg [31:0] z1775_assgn1775;
    reg [31:0] m3_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] m0_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5665_assgn5665;
    reg [31:0] z5665_assgn56650;
    reg [31:0] z5665_assgn56651;
    reg [31:0] z5665_assgn56652;
    reg [31:0] z1779_assgn1779;
    wire [31:0] p4_comar0_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5671_assgn5671;
    reg [31:0] z5671_assgn56710;
    reg [31:0] z5671_assgn56711;
    reg [31:0] z5671_assgn56712;
    reg [31:0] z1783_assgn1783;
    wire [31:0] i1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5675_assgn5675;
    reg [31:0] z5675_assgn56750;
    reg [31:0] z5675_assgn56751;
    reg [31:0] z5675_assgn56752;
    reg [31:0] z5675_assgn56753;
    reg [31:0] z5675_assgn56754;
    reg [31:0] z5675_assgn56755;
    reg [31:0] z1785_assgn1785;
    wire [31:0] i2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5679_assgn5679;
    reg [31:0] z5679_assgn56790;
    reg [31:0] z5679_assgn56791;
    reg [31:0] z5679_assgn56792;
    reg [31:0] z5679_assgn56793;
    reg [31:0] z5679_assgn56794;
    reg [31:0] z5679_assgn56795;
    reg [31:0] z1787_assgn1787;
    wire [31:0] i3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5683_assgn5683;
    reg [31:0] z5683_assgn56830;
    reg [31:0] z5683_assgn56831;
    reg [31:0] z5683_assgn56832;
    reg [31:0] z1790_assgn1790;
    reg [31:0] i2_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5687_assgn5687;
    reg [31:0] z5687_assgn56870;
    reg [31:0] z5687_assgn56871;
    reg [31:0] z5687_assgn56872;
    reg [31:0] z5687_assgn56873;
    reg [31:0] z5687_assgn56874;
    reg [31:0] z5687_assgn56875;
    reg [31:0] z1792_assgn1792;
    reg [31:0] i3_comar0_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] e0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] e1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r00_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m0_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5717_assgn5717;
    reg [31:0] z5717_assgn57170;
    reg [31:0] z5717_assgn57171;
    reg [31:0] z1819_assgn1819;
    wire [31:0] m1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5723_assgn5723;
    reg [31:0] z5723_assgn57230;
    reg [31:0] z5723_assgn57231;
    reg [31:0] z5723_assgn57232;
    reg [31:0] z5723_assgn57233;
    reg [31:0] z5723_assgn57234;
    reg [31:0] z1823_assgn1823;
    wire [31:0] m3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5727_assgn5727;
    reg [31:0] z5727_assgn57270;
    reg [31:0] z5727_assgn57271;
    reg [31:0] z5727_assgn57272;
    reg [31:0] z1826_assgn1826;
    reg [31:0] m1_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5731_assgn5731;
    reg [31:0] z5731_assgn57310;
    reg [31:0] z5731_assgn57311;
    reg [31:0] z5731_assgn57312;
    reg [31:0] z5731_assgn57313;
    reg [31:0] z5731_assgn57314;
    reg [31:0] z5731_assgn57315;
    reg [31:0] z1827_assgn1827;
    reg [31:0] m3_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] m0_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5737_assgn5737;
    reg [31:0] z5737_assgn57370;
    reg [31:0] z5737_assgn57371;
    reg [31:0] z5737_assgn57372;
    reg [31:0] z1831_assgn1831;
    wire [31:0] p4_comar1_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5743_assgn5743;
    reg [31:0] z5743_assgn57430;
    reg [31:0] z5743_assgn57431;
    reg [31:0] z5743_assgn57432;
    reg [31:0] z1835_assgn1835;
    wire [31:0] i1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5747_assgn5747;
    reg [31:0] z5747_assgn57470;
    reg [31:0] z5747_assgn57471;
    reg [31:0] z5747_assgn57472;
    reg [31:0] z5747_assgn57473;
    reg [31:0] z5747_assgn57474;
    reg [31:0] z5747_assgn57475;
    reg [31:0] z1837_assgn1837;
    wire [31:0] i2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5751_assgn5751;
    reg [31:0] z5751_assgn57510;
    reg [31:0] z5751_assgn57511;
    reg [31:0] z5751_assgn57512;
    reg [31:0] z5751_assgn57513;
    reg [31:0] z5751_assgn57514;
    reg [31:0] z5751_assgn57515;
    reg [31:0] z1839_assgn1839;
    wire [31:0] i3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5755_assgn5755;
    reg [31:0] z5755_assgn57550;
    reg [31:0] z5755_assgn57551;
    reg [31:0] z5755_assgn57552;
    reg [31:0] z1842_assgn1842;
    reg [31:0] i2_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5759_assgn5759;
    reg [31:0] z5759_assgn57590;
    reg [31:0] z5759_assgn57591;
    reg [31:0] z5759_assgn57592;
    reg [31:0] z5759_assgn57593;
    reg [31:0] z5759_assgn57594;
    reg [31:0] z5759_assgn57595;
    reg [31:0] z1844_assgn1844;
    reg [31:0] i3_comar1_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r00_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m0_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5793_assgn5793;
    reg [31:0] z5793_assgn57930;
    reg [31:0] z5793_assgn57931;
    reg [31:0] z1875_assgn1875;
    wire [31:0] m1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] m2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5799_assgn5799;
    reg [31:0] z5799_assgn57990;
    reg [31:0] z5799_assgn57991;
    reg [31:0] z5799_assgn57992;
    reg [31:0] z5799_assgn57993;
    reg [31:0] z5799_assgn57994;
    reg [31:0] z1879_assgn1879;
    wire [31:0] m3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5803_assgn5803;
    reg [31:0] z5803_assgn58030;
    reg [31:0] z5803_assgn58031;
    reg [31:0] z5803_assgn58032;
    reg [31:0] z1882_assgn1882;
    reg [31:0] m1_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5807_assgn5807;
    reg [31:0] z5807_assgn58070;
    reg [31:0] z5807_assgn58071;
    reg [31:0] z5807_assgn58072;
    reg [31:0] z5807_assgn58073;
    reg [31:0] z5807_assgn58074;
    reg [31:0] z5807_assgn58075;
    reg [31:0] z1883_assgn1883;
    reg [31:0] m3_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] m0_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    reg [31:0] m2_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5813_assgn5813;
    reg [31:0] z5813_assgn58130;
    reg [31:0] z5813_assgn58131;
    reg [31:0] z5813_assgn58132;
    reg [31:0] z1887_assgn1887;
    wire [31:0] p4_comar2_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5819_assgn5819;
    reg [31:0] z5819_assgn58190;
    reg [31:0] z5819_assgn58191;
    reg [31:0] z5819_assgn58192;
    reg [31:0] z1891_assgn1891;
    wire [31:0] i1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5823_assgn5823;
    reg [31:0] z5823_assgn58230;
    reg [31:0] z5823_assgn58231;
    reg [31:0] z5823_assgn58232;
    reg [31:0] z5823_assgn58233;
    reg [31:0] z5823_assgn58234;
    reg [31:0] z5823_assgn58235;
    reg [31:0] z1893_assgn1893;
    wire [31:0] i2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5827_assgn5827;
    reg [31:0] z5827_assgn58270;
    reg [31:0] z5827_assgn58271;
    reg [31:0] z5827_assgn58272;
    reg [31:0] z5827_assgn58273;
    reg [31:0] z5827_assgn58274;
    reg [31:0] z5827_assgn58275;
    reg [31:0] z1895_assgn1895;
    wire [31:0] i3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5831_assgn5831;
    reg [31:0] z5831_assgn58310;
    reg [31:0] z5831_assgn58311;
    reg [31:0] z5831_assgn58312;
    reg [31:0] z1898_assgn1898;
    reg [31:0] i2_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5835_assgn5835;
    reg [31:0] z5835_assgn58350;
    reg [31:0] z5835_assgn58351;
    reg [31:0] z5835_assgn58352;
    reg [31:0] z5835_assgn58353;
    reg [31:0] z5835_assgn58354;
    reg [31:0] z5835_assgn58355;
    reg [31:0] z1900_assgn1900;
    reg [31:0] i3_comar2_G4_mul5_G16_inv0_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0;
    reg [31:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] z5857_assgn5857;
    reg [31:0] z5857_assgn58570;
    reg [31:0] z5857_assgn58571;
    reg [31:0] z5857_assgn58572;
    reg [31:0] z5857_assgn58573;
    reg [31:0] z5857_assgn58574;
    reg [31:0] z5857_assgn58575;
    reg [31:0] z5857_assgn58576;
    reg [31:0] z5857_assgn58577;
    reg [31:0] z1919_assgn1919;
    wire [31:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [31:0] q0_G16_inv0_G256_inv0;
    wire [31:0] q1_G16_inv0_G256_inv0;
    wire [31:0] p0ls2_G16_inv0_G256_inv0;
    wire [31:0] z5867_assgn5867;
    reg [31:0] z5867_assgn58670;
    reg [31:0] z5867_assgn58671;
    reg [31:0] z5867_assgn58672;
    reg [31:0] z5867_assgn58673;
    reg [31:0] z5867_assgn58674;
    reg [31:0] z5867_assgn58675;
    reg [31:0] z5867_assgn58676;
    reg [31:0] z5867_assgn58677;
    reg [31:0] z1927_assgn1927;
    wire [31:0] p1ls2_G16_inv0_G256_inv0;
    wire [31:0] e0_G256_inv0;
    wire [31:0] e1_G256_inv0;
    wire [31:0] r00_G16_mul1_G256_inv0;
    wire [31:0] r10_G16_mul1_G256_inv0;
    wire [31:0] r20_G16_mul1_G256_inv0;
    wire [31:0] r30_G16_mul1_G256_inv0;
    wire [31:0] r40_G16_mul1_G256_inv0;
    wire [31:0] r50_G16_mul1_G256_inv0;
    wire [31:0] a0_0_G16_mul1_G256_inv0;
    wire [31:0] z5889_assgn5889;
    reg [31:0] z5889_assgn58890;
    reg [31:0] z5889_assgn58891;
    reg [31:0] z5889_assgn58892;
    reg [31:0] z5889_assgn58893;
    reg [31:0] z5889_assgn58894;
    reg [31:0] z5889_assgn58895;
    reg [31:0] z5889_assgn58896;
    reg [31:0] z5889_assgn58897;
    reg [31:0] z1947_assgn1947;
    wire [31:0] a1_0_G16_mul1_G256_inv0;
    wire [31:0] a0_G16_mul1_G256_inv0;
    wire [31:0] z5895_assgn5895;
    reg [31:0] z5895_assgn58950;
    reg [31:0] z5895_assgn58951;
    reg [31:0] z5895_assgn58952;
    reg [31:0] z5895_assgn58953;
    reg [31:0] z5895_assgn58954;
    reg [31:0] z5895_assgn58955;
    reg [31:0] z5895_assgn58956;
    reg [31:0] z5895_assgn58957;
    reg [31:0] z1951_assgn1951;
    wire [31:0] a1_G16_mul1_G256_inv0;
    wire [31:0] b0_G16_mul1_G256_inv0;
    wire [31:0] z5901_assgn5901;
    reg [31:0] z5901_assgn59010;
    reg [31:0] z5901_assgn59011;
    reg [31:0] z5901_assgn59012;
    reg [31:0] z5901_assgn59013;
    reg [31:0] z5901_assgn59014;
    reg [31:0] z5901_assgn59015;
    reg [31:0] z5901_assgn59016;
    reg [31:0] z5901_assgn59017;
    reg [31:0] z1955_assgn1955;
    wire [31:0] b1_G16_mul1_G256_inv0;
    wire [31:0] c0_0_G16_mul1_G256_inv0;
    wire [31:0] c1_0_G16_mul1_G256_inv0;
    wire [31:0] c0_G16_mul1_G256_inv0;
    wire [31:0] c1_G16_mul1_G256_inv0;
    wire [31:0] d0_G16_mul1_G256_inv0;
    wire [31:0] d1_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G16_mul1_G256_inv0;
    wire [31:0] cxord_0_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G16_mul1_G256_inv0;
    wire [31:0] cxord_1_G16_mul1_G256_inv0;
    wire [31:0] r00_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r10_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r20_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r30_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r40_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r50_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5939_assgn5939;
    reg [31:0] z5939_assgn59390;
    reg [31:0] z5939_assgn59391;
    reg [31:0] z5939_assgn59392;
    reg [31:0] z5939_assgn59393;
    reg [31:0] z5939_assgn59394;
    reg [31:0] z5939_assgn59395;
    reg [31:0] z5939_assgn59396;
    reg [31:0] z5939_assgn59397;
    reg [31:0] z1991_assgn1991;
    wire [31:0] a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5945_assgn5945;
    reg [31:0] z5945_assgn59450;
    reg [31:0] z5945_assgn59451;
    reg [31:0] z5945_assgn59452;
    reg [31:0] z5945_assgn59453;
    reg [31:0] z5945_assgn59454;
    reg [31:0] z5945_assgn59455;
    reg [31:0] z5945_assgn59456;
    reg [31:0] z5945_assgn59457;
    reg [31:0] z1995_assgn1995;
    wire [31:0] a1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5951_assgn5951;
    reg [31:0] z5951_assgn59510;
    reg [31:0] z5951_assgn59511;
    reg [31:0] z5951_assgn59512;
    reg [31:0] z5951_assgn59513;
    reg [31:0] z5951_assgn59514;
    reg [31:0] z5951_assgn59515;
    reg [31:0] z5951_assgn59516;
    reg [31:0] z5951_assgn59517;
    reg [31:0] z1999_assgn1999;
    wire [31:0] b1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] c1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] d1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r00_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m0_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5993_assgn5993;
    reg [31:0] z5993_assgn59930;
    reg [31:0] z5993_assgn59931;
    reg [31:0] z5993_assgn59932;
    reg [31:0] z5993_assgn59933;
    reg [31:0] z5993_assgn59934;
    reg [31:0] z5993_assgn59935;
    reg [31:0] z5993_assgn59936;
    reg [31:0] z5993_assgn59937;
    reg [31:0] z2039_assgn2039;
    wire [31:0] m3_comar0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m0_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z5999_assgn5999;
    reg [31:0] z5999_assgn59990;
    reg [31:0] z5999_assgn59991;
    reg [31:0] z5999_assgn59992;
    reg [31:0] z5999_assgn59993;
    reg [31:0] z5999_assgn59994;
    reg [31:0] z5999_assgn59995;
    reg [31:0] z5999_assgn59996;
    reg [31:0] z5999_assgn59997;
    reg [31:0] z5999_assgn59998;
    reg [31:0] z2043_assgn2043;
    reg [31:0] m3_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m2_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6005_assgn6005;
    reg [31:0] z6005_assgn60050;
    reg [31:0] z6005_assgn60051;
    reg [31:0] z6005_assgn60052;
    reg [31:0] z6005_assgn60053;
    reg [31:0] z6005_assgn60054;
    reg [31:0] z6005_assgn60055;
    reg [31:0] z6005_assgn60056;
    reg [31:0] z6005_assgn60057;
    reg [31:0] z6005_assgn60058;
    reg [31:0] z2047_assgn2047;
    wire [31:0] p4_comar0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6013_assgn6013;
    reg [31:0] z6013_assgn60130;
    reg [31:0] z6013_assgn60131;
    reg [31:0] z6013_assgn60132;
    reg [31:0] z6013_assgn60133;
    reg [31:0] z6013_assgn60134;
    reg [31:0] z6013_assgn60135;
    reg [31:0] z6013_assgn60136;
    reg [31:0] z6013_assgn60137;
    reg [31:0] z6013_assgn60138;
    reg [31:0] z2053_assgn2053;
    wire [31:0] i2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6017_assgn6017;
    reg [31:0] z6017_assgn60170;
    reg [31:0] z6017_assgn60171;
    reg [31:0] z6017_assgn60172;
    reg [31:0] z6017_assgn60173;
    reg [31:0] z6017_assgn60174;
    reg [31:0] z6017_assgn60175;
    reg [31:0] z6017_assgn60176;
    reg [31:0] z6017_assgn60177;
    reg [31:0] z6017_assgn60178;
    reg [31:0] z2055_assgn2055;
    wire [31:0] i3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6021_assgn6021;
    reg [31:0] z6021_assgn60210;
    reg [31:0] z6021_assgn60211;
    reg [31:0] z6021_assgn60212;
    reg [31:0] z6021_assgn60213;
    reg [31:0] z6021_assgn60214;
    reg [31:0] z6021_assgn60215;
    reg [31:0] z6021_assgn60216;
    reg [31:0] z6021_assgn60217;
    reg [31:0] z6021_assgn60218;
    reg [31:0] z2058_assgn2058;
    reg [31:0] i2_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6025_assgn6025;
    reg [31:0] z6025_assgn60250;
    reg [31:0] z6025_assgn60251;
    reg [31:0] z6025_assgn60252;
    reg [31:0] z6025_assgn60253;
    reg [31:0] z6025_assgn60254;
    reg [31:0] z6025_assgn60255;
    reg [31:0] z6025_assgn60256;
    reg [31:0] z6025_assgn60257;
    reg [31:0] z6025_assgn60258;
    reg [31:0] z2060_assgn2060;
    reg [31:0] i3_comar0_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] e0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] e1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r00_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m0_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6059_assgn6059;
    reg [31:0] z6059_assgn60590;
    reg [31:0] z6059_assgn60591;
    reg [31:0] z6059_assgn60592;
    reg [31:0] z6059_assgn60593;
    reg [31:0] z6059_assgn60594;
    reg [31:0] z6059_assgn60595;
    reg [31:0] z6059_assgn60596;
    reg [31:0] z6059_assgn60597;
    reg [31:0] z2091_assgn2091;
    wire [31:0] m3_comar1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m0_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6065_assgn6065;
    reg [31:0] z6065_assgn60650;
    reg [31:0] z6065_assgn60651;
    reg [31:0] z6065_assgn60652;
    reg [31:0] z6065_assgn60653;
    reg [31:0] z6065_assgn60654;
    reg [31:0] z6065_assgn60655;
    reg [31:0] z6065_assgn60656;
    reg [31:0] z6065_assgn60657;
    reg [31:0] z6065_assgn60658;
    reg [31:0] z2095_assgn2095;
    reg [31:0] m3_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m2_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6071_assgn6071;
    reg [31:0] z6071_assgn60710;
    reg [31:0] z6071_assgn60711;
    reg [31:0] z6071_assgn60712;
    reg [31:0] z6071_assgn60713;
    reg [31:0] z6071_assgn60714;
    reg [31:0] z6071_assgn60715;
    reg [31:0] z6071_assgn60716;
    reg [31:0] z6071_assgn60717;
    reg [31:0] z6071_assgn60718;
    reg [31:0] z2099_assgn2099;
    wire [31:0] p4_comar1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6079_assgn6079;
    reg [31:0] z6079_assgn60790;
    reg [31:0] z6079_assgn60791;
    reg [31:0] z6079_assgn60792;
    reg [31:0] z6079_assgn60793;
    reg [31:0] z6079_assgn60794;
    reg [31:0] z6079_assgn60795;
    reg [31:0] z6079_assgn60796;
    reg [31:0] z6079_assgn60797;
    reg [31:0] z6079_assgn60798;
    reg [31:0] z2105_assgn2105;
    wire [31:0] i2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6083_assgn6083;
    reg [31:0] z6083_assgn60830;
    reg [31:0] z6083_assgn60831;
    reg [31:0] z6083_assgn60832;
    reg [31:0] z6083_assgn60833;
    reg [31:0] z6083_assgn60834;
    reg [31:0] z6083_assgn60835;
    reg [31:0] z6083_assgn60836;
    reg [31:0] z6083_assgn60837;
    reg [31:0] z6083_assgn60838;
    reg [31:0] z2107_assgn2107;
    wire [31:0] i3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6087_assgn6087;
    reg [31:0] z6087_assgn60870;
    reg [31:0] z6087_assgn60871;
    reg [31:0] z6087_assgn60872;
    reg [31:0] z6087_assgn60873;
    reg [31:0] z6087_assgn60874;
    reg [31:0] z6087_assgn60875;
    reg [31:0] z6087_assgn60876;
    reg [31:0] z6087_assgn60877;
    reg [31:0] z6087_assgn60878;
    reg [31:0] z2110_assgn2110;
    reg [31:0] i2_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6091_assgn6091;
    reg [31:0] z6091_assgn60910;
    reg [31:0] z6091_assgn60911;
    reg [31:0] z6091_assgn60912;
    reg [31:0] z6091_assgn60913;
    reg [31:0] z6091_assgn60914;
    reg [31:0] z6091_assgn60915;
    reg [31:0] z6091_assgn60916;
    reg [31:0] z6091_assgn60917;
    reg [31:0] z6091_assgn60918;
    reg [31:0] z2112_assgn2112;
    reg [31:0] i3_comar1_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r00_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m0_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] m2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6129_assgn6129;
    reg [31:0] z6129_assgn61290;
    reg [31:0] z6129_assgn61291;
    reg [31:0] z6129_assgn61292;
    reg [31:0] z6129_assgn61293;
    reg [31:0] z6129_assgn61294;
    reg [31:0] z6129_assgn61295;
    reg [31:0] z6129_assgn61296;
    reg [31:0] z6129_assgn61297;
    reg [31:0] z2147_assgn2147;
    wire [31:0] m3_comar2_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m0_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6135_assgn6135;
    reg [31:0] z6135_assgn61350;
    reg [31:0] z6135_assgn61351;
    reg [31:0] z6135_assgn61352;
    reg [31:0] z6135_assgn61353;
    reg [31:0] z6135_assgn61354;
    reg [31:0] z6135_assgn61355;
    reg [31:0] z6135_assgn61356;
    reg [31:0] z6135_assgn61357;
    reg [31:0] z6135_assgn61358;
    reg [31:0] z2151_assgn2151;
    reg [31:0] m3_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] m2_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6141_assgn6141;
    reg [31:0] z6141_assgn61410;
    reg [31:0] z6141_assgn61411;
    reg [31:0] z6141_assgn61412;
    reg [31:0] z6141_assgn61413;
    reg [31:0] z6141_assgn61414;
    reg [31:0] z6141_assgn61415;
    reg [31:0] z6141_assgn61416;
    reg [31:0] z6141_assgn61417;
    reg [31:0] z6141_assgn61418;
    reg [31:0] z2155_assgn2155;
    wire [31:0] p4_comar2_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6149_assgn6149;
    reg [31:0] z6149_assgn61490;
    reg [31:0] z6149_assgn61491;
    reg [31:0] z6149_assgn61492;
    reg [31:0] z6149_assgn61493;
    reg [31:0] z6149_assgn61494;
    reg [31:0] z6149_assgn61495;
    reg [31:0] z6149_assgn61496;
    reg [31:0] z6149_assgn61497;
    reg [31:0] z6149_assgn61498;
    reg [31:0] z2161_assgn2161;
    wire [31:0] i2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6153_assgn6153;
    reg [31:0] z6153_assgn61530;
    reg [31:0] z6153_assgn61531;
    reg [31:0] z6153_assgn61532;
    reg [31:0] z6153_assgn61533;
    reg [31:0] z6153_assgn61534;
    reg [31:0] z6153_assgn61535;
    reg [31:0] z6153_assgn61536;
    reg [31:0] z6153_assgn61537;
    reg [31:0] z6153_assgn61538;
    reg [31:0] z2163_assgn2163;
    wire [31:0] i3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6157_assgn6157;
    reg [31:0] z6157_assgn61570;
    reg [31:0] z6157_assgn61571;
    reg [31:0] z6157_assgn61572;
    reg [31:0] z6157_assgn61573;
    reg [31:0] z6157_assgn61574;
    reg [31:0] z6157_assgn61575;
    reg [31:0] z6157_assgn61576;
    reg [31:0] z6157_assgn61577;
    reg [31:0] z6157_assgn61578;
    reg [31:0] z2166_assgn2166;
    reg [31:0] i2_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6161_assgn6161;
    reg [31:0] z6161_assgn61610;
    reg [31:0] z6161_assgn61611;
    reg [31:0] z6161_assgn61612;
    reg [31:0] z6161_assgn61613;
    reg [31:0] z6161_assgn61614;
    reg [31:0] z6161_assgn61615;
    reg [31:0] z6161_assgn61616;
    reg [31:0] z6161_assgn61617;
    reg [31:0] z6161_assgn61618;
    reg [31:0] z2168_assgn2168;
    reg [31:0] i3_comar2_G4_mul0_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0;
    reg [31:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] z6183_assgn6183;
    reg [31:0] z6183_assgn61830;
    reg [31:0] z6183_assgn61831;
    reg [31:0] z6183_assgn61832;
    reg [31:0] z6183_assgn61833;
    reg [31:0] z6183_assgn61834;
    reg [31:0] z6183_assgn61835;
    reg [31:0] z6183_assgn61836;
    reg [31:0] z6183_assgn61837;
    reg [31:0] z6183_assgn61838;
    reg [31:0] z6183_assgn61839;
    reg [31:0] z6183_assgn618310;
    reg [31:0] z2187_assgn2187;
    wire [31:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [31:0] e0_G16_mul1_G256_inv0;
    wire [31:0] e1_G16_mul1_G256_inv0;
    wire [31:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z6193_assgn6193;
    reg [31:0] z6193_assgn61930;
    reg [31:0] z6193_assgn61931;
    reg [31:0] z6193_assgn61932;
    reg [31:0] z6193_assgn61933;
    reg [31:0] z6193_assgn61934;
    reg [31:0] z6193_assgn61935;
    reg [31:0] z6193_assgn61936;
    reg [31:0] z6193_assgn61937;
    reg [31:0] z6193_assgn61938;
    reg [31:0] z6193_assgn61939;
    reg [31:0] z6193_assgn619310;
    reg [31:0] z2195_assgn2195;
    wire [31:0] a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z6199_assgn6199;
    reg [31:0] z6199_assgn61990;
    reg [31:0] z6199_assgn61991;
    reg [31:0] z6199_assgn61992;
    reg [31:0] z6199_assgn61993;
    reg [31:0] z6199_assgn61994;
    reg [31:0] z6199_assgn61995;
    reg [31:0] z6199_assgn61996;
    reg [31:0] z6199_assgn61997;
    reg [31:0] z6199_assgn61998;
    reg [31:0] z6199_assgn61999;
    reg [31:0] z6199_assgn619910;
    reg [31:0] z2199_assgn2199;
    wire [31:0] a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z6205_assgn6205;
    reg [31:0] z6205_assgn62050;
    reg [31:0] z6205_assgn62051;
    reg [31:0] z6205_assgn62052;
    reg [31:0] z6205_assgn62053;
    reg [31:0] z6205_assgn62054;
    reg [31:0] z6205_assgn62055;
    reg [31:0] z6205_assgn62056;
    reg [31:0] z6205_assgn62057;
    reg [31:0] z6205_assgn62058;
    reg [31:0] z6205_assgn62059;
    reg [31:0] z6205_assgn620510;
    reg [31:0] z2203_assgn2203;
    wire [31:0] b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] z6217_assgn6217;
    reg [31:0] z6217_assgn62170;
    reg [31:0] z6217_assgn62171;
    reg [31:0] z6217_assgn62172;
    reg [31:0] z6217_assgn62173;
    reg [31:0] z6217_assgn62174;
    reg [31:0] z6217_assgn62175;
    reg [31:0] z6217_assgn62176;
    reg [31:0] z6217_assgn62177;
    reg [31:0] z6217_assgn62178;
    reg [31:0] z6217_assgn62179;
    reg [31:0] z6217_assgn621710;
    reg [31:0] z2213_assgn2213;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [31:0] e01_G16_mul1_G256_inv0;
    wire [31:0] e11_G16_mul1_G256_inv0;
    wire [31:0] r00_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r10_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r20_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r30_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r40_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r50_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6241_assgn6241;
    reg [31:0] z6241_assgn62410;
    reg [31:0] z6241_assgn62411;
    reg [31:0] z6241_assgn62412;
    reg [31:0] z6241_assgn62413;
    reg [31:0] z6241_assgn62414;
    reg [31:0] z6241_assgn62415;
    reg [31:0] z6241_assgn62416;
    reg [31:0] z6241_assgn62417;
    reg [31:0] z2235_assgn2235;
    wire [31:0] a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6247_assgn6247;
    reg [31:0] z6247_assgn62470;
    reg [31:0] z6247_assgn62471;
    reg [31:0] z6247_assgn62472;
    reg [31:0] z6247_assgn62473;
    reg [31:0] z6247_assgn62474;
    reg [31:0] z6247_assgn62475;
    reg [31:0] z6247_assgn62476;
    reg [31:0] z6247_assgn62477;
    reg [31:0] z2239_assgn2239;
    wire [31:0] a1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6253_assgn6253;
    reg [31:0] z6253_assgn62530;
    reg [31:0] z6253_assgn62531;
    reg [31:0] z6253_assgn62532;
    reg [31:0] z6253_assgn62533;
    reg [31:0] z6253_assgn62534;
    reg [31:0] z6253_assgn62535;
    reg [31:0] z6253_assgn62536;
    reg [31:0] z6253_assgn62537;
    reg [31:0] z2243_assgn2243;
    wire [31:0] b1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] c1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] d1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r00_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m0_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6295_assgn6295;
    reg [31:0] z6295_assgn62950;
    reg [31:0] z6295_assgn62951;
    reg [31:0] z6295_assgn62952;
    reg [31:0] z6295_assgn62953;
    reg [31:0] z6295_assgn62954;
    reg [31:0] z6295_assgn62955;
    reg [31:0] z6295_assgn62956;
    reg [31:0] z6295_assgn62957;
    reg [31:0] z2283_assgn2283;
    wire [31:0] m3_comar0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m0_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6301_assgn6301;
    reg [31:0] z6301_assgn63010;
    reg [31:0] z6301_assgn63011;
    reg [31:0] z6301_assgn63012;
    reg [31:0] z6301_assgn63013;
    reg [31:0] z6301_assgn63014;
    reg [31:0] z6301_assgn63015;
    reg [31:0] z6301_assgn63016;
    reg [31:0] z6301_assgn63017;
    reg [31:0] z6301_assgn63018;
    reg [31:0] z2287_assgn2287;
    reg [31:0] m3_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m2_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6307_assgn6307;
    reg [31:0] z6307_assgn63070;
    reg [31:0] z6307_assgn63071;
    reg [31:0] z6307_assgn63072;
    reg [31:0] z6307_assgn63073;
    reg [31:0] z6307_assgn63074;
    reg [31:0] z6307_assgn63075;
    reg [31:0] z6307_assgn63076;
    reg [31:0] z6307_assgn63077;
    reg [31:0] z6307_assgn63078;
    reg [31:0] z2291_assgn2291;
    wire [31:0] p4_comar0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6315_assgn6315;
    reg [31:0] z6315_assgn63150;
    reg [31:0] z6315_assgn63151;
    reg [31:0] z6315_assgn63152;
    reg [31:0] z6315_assgn63153;
    reg [31:0] z6315_assgn63154;
    reg [31:0] z6315_assgn63155;
    reg [31:0] z6315_assgn63156;
    reg [31:0] z6315_assgn63157;
    reg [31:0] z6315_assgn63158;
    reg [31:0] z2297_assgn2297;
    wire [31:0] i2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6319_assgn6319;
    reg [31:0] z6319_assgn63190;
    reg [31:0] z6319_assgn63191;
    reg [31:0] z6319_assgn63192;
    reg [31:0] z6319_assgn63193;
    reg [31:0] z6319_assgn63194;
    reg [31:0] z6319_assgn63195;
    reg [31:0] z6319_assgn63196;
    reg [31:0] z6319_assgn63197;
    reg [31:0] z6319_assgn63198;
    reg [31:0] z2299_assgn2299;
    wire [31:0] i3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6323_assgn6323;
    reg [31:0] z6323_assgn63230;
    reg [31:0] z6323_assgn63231;
    reg [31:0] z6323_assgn63232;
    reg [31:0] z6323_assgn63233;
    reg [31:0] z6323_assgn63234;
    reg [31:0] z6323_assgn63235;
    reg [31:0] z6323_assgn63236;
    reg [31:0] z6323_assgn63237;
    reg [31:0] z6323_assgn63238;
    reg [31:0] z2302_assgn2302;
    reg [31:0] i2_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6327_assgn6327;
    reg [31:0] z6327_assgn63270;
    reg [31:0] z6327_assgn63271;
    reg [31:0] z6327_assgn63272;
    reg [31:0] z6327_assgn63273;
    reg [31:0] z6327_assgn63274;
    reg [31:0] z6327_assgn63275;
    reg [31:0] z6327_assgn63276;
    reg [31:0] z6327_assgn63277;
    reg [31:0] z6327_assgn63278;
    reg [31:0] z2304_assgn2304;
    reg [31:0] i3_comar0_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] e0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] e1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r00_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m0_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6361_assgn6361;
    reg [31:0] z6361_assgn63610;
    reg [31:0] z6361_assgn63611;
    reg [31:0] z6361_assgn63612;
    reg [31:0] z6361_assgn63613;
    reg [31:0] z6361_assgn63614;
    reg [31:0] z6361_assgn63615;
    reg [31:0] z6361_assgn63616;
    reg [31:0] z6361_assgn63617;
    reg [31:0] z2335_assgn2335;
    wire [31:0] m3_comar1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m0_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6367_assgn6367;
    reg [31:0] z6367_assgn63670;
    reg [31:0] z6367_assgn63671;
    reg [31:0] z6367_assgn63672;
    reg [31:0] z6367_assgn63673;
    reg [31:0] z6367_assgn63674;
    reg [31:0] z6367_assgn63675;
    reg [31:0] z6367_assgn63676;
    reg [31:0] z6367_assgn63677;
    reg [31:0] z6367_assgn63678;
    reg [31:0] z2339_assgn2339;
    reg [31:0] m3_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m2_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6373_assgn6373;
    reg [31:0] z6373_assgn63730;
    reg [31:0] z6373_assgn63731;
    reg [31:0] z6373_assgn63732;
    reg [31:0] z6373_assgn63733;
    reg [31:0] z6373_assgn63734;
    reg [31:0] z6373_assgn63735;
    reg [31:0] z6373_assgn63736;
    reg [31:0] z6373_assgn63737;
    reg [31:0] z6373_assgn63738;
    reg [31:0] z2343_assgn2343;
    wire [31:0] p4_comar1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6381_assgn6381;
    reg [31:0] z6381_assgn63810;
    reg [31:0] z6381_assgn63811;
    reg [31:0] z6381_assgn63812;
    reg [31:0] z6381_assgn63813;
    reg [31:0] z6381_assgn63814;
    reg [31:0] z6381_assgn63815;
    reg [31:0] z6381_assgn63816;
    reg [31:0] z6381_assgn63817;
    reg [31:0] z6381_assgn63818;
    reg [31:0] z2349_assgn2349;
    wire [31:0] i2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6385_assgn6385;
    reg [31:0] z6385_assgn63850;
    reg [31:0] z6385_assgn63851;
    reg [31:0] z6385_assgn63852;
    reg [31:0] z6385_assgn63853;
    reg [31:0] z6385_assgn63854;
    reg [31:0] z6385_assgn63855;
    reg [31:0] z6385_assgn63856;
    reg [31:0] z6385_assgn63857;
    reg [31:0] z6385_assgn63858;
    reg [31:0] z2351_assgn2351;
    wire [31:0] i3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6389_assgn6389;
    reg [31:0] z6389_assgn63890;
    reg [31:0] z6389_assgn63891;
    reg [31:0] z6389_assgn63892;
    reg [31:0] z6389_assgn63893;
    reg [31:0] z6389_assgn63894;
    reg [31:0] z6389_assgn63895;
    reg [31:0] z6389_assgn63896;
    reg [31:0] z6389_assgn63897;
    reg [31:0] z6389_assgn63898;
    reg [31:0] z2354_assgn2354;
    reg [31:0] i2_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6393_assgn6393;
    reg [31:0] z6393_assgn63930;
    reg [31:0] z6393_assgn63931;
    reg [31:0] z6393_assgn63932;
    reg [31:0] z6393_assgn63933;
    reg [31:0] z6393_assgn63934;
    reg [31:0] z6393_assgn63935;
    reg [31:0] z6393_assgn63936;
    reg [31:0] z6393_assgn63937;
    reg [31:0] z6393_assgn63938;
    reg [31:0] z2356_assgn2356;
    reg [31:0] i3_comar1_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r00_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m0_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] m2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6431_assgn6431;
    reg [31:0] z6431_assgn64310;
    reg [31:0] z6431_assgn64311;
    reg [31:0] z6431_assgn64312;
    reg [31:0] z6431_assgn64313;
    reg [31:0] z6431_assgn64314;
    reg [31:0] z6431_assgn64315;
    reg [31:0] z6431_assgn64316;
    reg [31:0] z6431_assgn64317;
    reg [31:0] z2391_assgn2391;
    wire [31:0] m3_comar2_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m0_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6437_assgn6437;
    reg [31:0] z6437_assgn64370;
    reg [31:0] z6437_assgn64371;
    reg [31:0] z6437_assgn64372;
    reg [31:0] z6437_assgn64373;
    reg [31:0] z6437_assgn64374;
    reg [31:0] z6437_assgn64375;
    reg [31:0] z6437_assgn64376;
    reg [31:0] z6437_assgn64377;
    reg [31:0] z6437_assgn64378;
    reg [31:0] z2395_assgn2395;
    reg [31:0] m3_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] m2_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6443_assgn6443;
    reg [31:0] z6443_assgn64430;
    reg [31:0] z6443_assgn64431;
    reg [31:0] z6443_assgn64432;
    reg [31:0] z6443_assgn64433;
    reg [31:0] z6443_assgn64434;
    reg [31:0] z6443_assgn64435;
    reg [31:0] z6443_assgn64436;
    reg [31:0] z6443_assgn64437;
    reg [31:0] z6443_assgn64438;
    reg [31:0] z2399_assgn2399;
    wire [31:0] p4_comar2_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6451_assgn6451;
    reg [31:0] z6451_assgn64510;
    reg [31:0] z6451_assgn64511;
    reg [31:0] z6451_assgn64512;
    reg [31:0] z6451_assgn64513;
    reg [31:0] z6451_assgn64514;
    reg [31:0] z6451_assgn64515;
    reg [31:0] z6451_assgn64516;
    reg [31:0] z6451_assgn64517;
    reg [31:0] z6451_assgn64518;
    reg [31:0] z2405_assgn2405;
    wire [31:0] i2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6455_assgn6455;
    reg [31:0] z6455_assgn64550;
    reg [31:0] z6455_assgn64551;
    reg [31:0] z6455_assgn64552;
    reg [31:0] z6455_assgn64553;
    reg [31:0] z6455_assgn64554;
    reg [31:0] z6455_assgn64555;
    reg [31:0] z6455_assgn64556;
    reg [31:0] z6455_assgn64557;
    reg [31:0] z6455_assgn64558;
    reg [31:0] z2407_assgn2407;
    wire [31:0] i3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6459_assgn6459;
    reg [31:0] z6459_assgn64590;
    reg [31:0] z6459_assgn64591;
    reg [31:0] z6459_assgn64592;
    reg [31:0] z6459_assgn64593;
    reg [31:0] z6459_assgn64594;
    reg [31:0] z6459_assgn64595;
    reg [31:0] z6459_assgn64596;
    reg [31:0] z6459_assgn64597;
    reg [31:0] z6459_assgn64598;
    reg [31:0] z2410_assgn2410;
    reg [31:0] i2_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6463_assgn6463;
    reg [31:0] z6463_assgn64630;
    reg [31:0] z6463_assgn64631;
    reg [31:0] z6463_assgn64632;
    reg [31:0] z6463_assgn64633;
    reg [31:0] z6463_assgn64634;
    reg [31:0] z6463_assgn64635;
    reg [31:0] z6463_assgn64636;
    reg [31:0] z6463_assgn64637;
    reg [31:0] z6463_assgn64638;
    reg [31:0] z2412_assgn2412;
    reg [31:0] i3_comar2_G4_mul1_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0;
    reg [31:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] z6485_assgn6485;
    reg [31:0] z6485_assgn64850;
    reg [31:0] z6485_assgn64851;
    reg [31:0] z6485_assgn64852;
    reg [31:0] z6485_assgn64853;
    reg [31:0] z6485_assgn64854;
    reg [31:0] z6485_assgn64855;
    reg [31:0] z6485_assgn64856;
    reg [31:0] z6485_assgn64857;
    reg [31:0] z6485_assgn64858;
    reg [31:0] z6485_assgn64859;
    reg [31:0] z6485_assgn648510;
    reg [31:0] z2431_assgn2431;
    wire [31:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [31:0] p0_0_G16_mul1_G256_inv0;
    wire [31:0] p1_0_G16_mul1_G256_inv0;
    wire [31:0] p0_G16_mul1_G256_inv0;
    wire [31:0] p1_G16_mul1_G256_inv0;
    wire [31:0] r00_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r10_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r20_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r30_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r40_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r50_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6511_assgn6511;
    reg [31:0] z6511_assgn65110;
    reg [31:0] z6511_assgn65111;
    reg [31:0] z6511_assgn65112;
    reg [31:0] z6511_assgn65113;
    reg [31:0] z6511_assgn65114;
    reg [31:0] z6511_assgn65115;
    reg [31:0] z6511_assgn65116;
    reg [31:0] z6511_assgn65117;
    reg [31:0] z2455_assgn2455;
    wire [31:0] a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6517_assgn6517;
    reg [31:0] z6517_assgn65170;
    reg [31:0] z6517_assgn65171;
    reg [31:0] z6517_assgn65172;
    reg [31:0] z6517_assgn65173;
    reg [31:0] z6517_assgn65174;
    reg [31:0] z6517_assgn65175;
    reg [31:0] z6517_assgn65176;
    reg [31:0] z6517_assgn65177;
    reg [31:0] z2459_assgn2459;
    wire [31:0] a1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6523_assgn6523;
    reg [31:0] z6523_assgn65230;
    reg [31:0] z6523_assgn65231;
    reg [31:0] z6523_assgn65232;
    reg [31:0] z6523_assgn65233;
    reg [31:0] z6523_assgn65234;
    reg [31:0] z6523_assgn65235;
    reg [31:0] z6523_assgn65236;
    reg [31:0] z6523_assgn65237;
    reg [31:0] z2463_assgn2463;
    wire [31:0] b1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] c1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] d1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r00_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m0_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6565_assgn6565;
    reg [31:0] z6565_assgn65650;
    reg [31:0] z6565_assgn65651;
    reg [31:0] z6565_assgn65652;
    reg [31:0] z6565_assgn65653;
    reg [31:0] z6565_assgn65654;
    reg [31:0] z6565_assgn65655;
    reg [31:0] z6565_assgn65656;
    reg [31:0] z6565_assgn65657;
    reg [31:0] z2503_assgn2503;
    wire [31:0] m3_comar0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m0_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6571_assgn6571;
    reg [31:0] z6571_assgn65710;
    reg [31:0] z6571_assgn65711;
    reg [31:0] z6571_assgn65712;
    reg [31:0] z6571_assgn65713;
    reg [31:0] z6571_assgn65714;
    reg [31:0] z6571_assgn65715;
    reg [31:0] z6571_assgn65716;
    reg [31:0] z6571_assgn65717;
    reg [31:0] z6571_assgn65718;
    reg [31:0] z2507_assgn2507;
    reg [31:0] m3_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m2_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6577_assgn6577;
    reg [31:0] z6577_assgn65770;
    reg [31:0] z6577_assgn65771;
    reg [31:0] z6577_assgn65772;
    reg [31:0] z6577_assgn65773;
    reg [31:0] z6577_assgn65774;
    reg [31:0] z6577_assgn65775;
    reg [31:0] z6577_assgn65776;
    reg [31:0] z6577_assgn65777;
    reg [31:0] z6577_assgn65778;
    reg [31:0] z2511_assgn2511;
    wire [31:0] p4_comar0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6585_assgn6585;
    reg [31:0] z6585_assgn65850;
    reg [31:0] z6585_assgn65851;
    reg [31:0] z6585_assgn65852;
    reg [31:0] z6585_assgn65853;
    reg [31:0] z6585_assgn65854;
    reg [31:0] z6585_assgn65855;
    reg [31:0] z6585_assgn65856;
    reg [31:0] z6585_assgn65857;
    reg [31:0] z6585_assgn65858;
    reg [31:0] z2517_assgn2517;
    wire [31:0] i2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6589_assgn6589;
    reg [31:0] z6589_assgn65890;
    reg [31:0] z6589_assgn65891;
    reg [31:0] z6589_assgn65892;
    reg [31:0] z6589_assgn65893;
    reg [31:0] z6589_assgn65894;
    reg [31:0] z6589_assgn65895;
    reg [31:0] z6589_assgn65896;
    reg [31:0] z6589_assgn65897;
    reg [31:0] z6589_assgn65898;
    reg [31:0] z2519_assgn2519;
    wire [31:0] i3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6593_assgn6593;
    reg [31:0] z6593_assgn65930;
    reg [31:0] z6593_assgn65931;
    reg [31:0] z6593_assgn65932;
    reg [31:0] z6593_assgn65933;
    reg [31:0] z6593_assgn65934;
    reg [31:0] z6593_assgn65935;
    reg [31:0] z6593_assgn65936;
    reg [31:0] z6593_assgn65937;
    reg [31:0] z6593_assgn65938;
    reg [31:0] z2522_assgn2522;
    reg [31:0] i2_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6597_assgn6597;
    reg [31:0] z6597_assgn65970;
    reg [31:0] z6597_assgn65971;
    reg [31:0] z6597_assgn65972;
    reg [31:0] z6597_assgn65973;
    reg [31:0] z6597_assgn65974;
    reg [31:0] z6597_assgn65975;
    reg [31:0] z6597_assgn65976;
    reg [31:0] z6597_assgn65977;
    reg [31:0] z6597_assgn65978;
    reg [31:0] z2524_assgn2524;
    reg [31:0] i3_comar0_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] e0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] e1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r00_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m0_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6631_assgn6631;
    reg [31:0] z6631_assgn66310;
    reg [31:0] z6631_assgn66311;
    reg [31:0] z6631_assgn66312;
    reg [31:0] z6631_assgn66313;
    reg [31:0] z6631_assgn66314;
    reg [31:0] z6631_assgn66315;
    reg [31:0] z6631_assgn66316;
    reg [31:0] z6631_assgn66317;
    reg [31:0] z2555_assgn2555;
    wire [31:0] m3_comar1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m0_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6637_assgn6637;
    reg [31:0] z6637_assgn66370;
    reg [31:0] z6637_assgn66371;
    reg [31:0] z6637_assgn66372;
    reg [31:0] z6637_assgn66373;
    reg [31:0] z6637_assgn66374;
    reg [31:0] z6637_assgn66375;
    reg [31:0] z6637_assgn66376;
    reg [31:0] z6637_assgn66377;
    reg [31:0] z6637_assgn66378;
    reg [31:0] z2559_assgn2559;
    reg [31:0] m3_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m2_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6643_assgn6643;
    reg [31:0] z6643_assgn66430;
    reg [31:0] z6643_assgn66431;
    reg [31:0] z6643_assgn66432;
    reg [31:0] z6643_assgn66433;
    reg [31:0] z6643_assgn66434;
    reg [31:0] z6643_assgn66435;
    reg [31:0] z6643_assgn66436;
    reg [31:0] z6643_assgn66437;
    reg [31:0] z6643_assgn66438;
    reg [31:0] z2563_assgn2563;
    wire [31:0] p4_comar1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6651_assgn6651;
    reg [31:0] z6651_assgn66510;
    reg [31:0] z6651_assgn66511;
    reg [31:0] z6651_assgn66512;
    reg [31:0] z6651_assgn66513;
    reg [31:0] z6651_assgn66514;
    reg [31:0] z6651_assgn66515;
    reg [31:0] z6651_assgn66516;
    reg [31:0] z6651_assgn66517;
    reg [31:0] z6651_assgn66518;
    reg [31:0] z2569_assgn2569;
    wire [31:0] i2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6655_assgn6655;
    reg [31:0] z6655_assgn66550;
    reg [31:0] z6655_assgn66551;
    reg [31:0] z6655_assgn66552;
    reg [31:0] z6655_assgn66553;
    reg [31:0] z6655_assgn66554;
    reg [31:0] z6655_assgn66555;
    reg [31:0] z6655_assgn66556;
    reg [31:0] z6655_assgn66557;
    reg [31:0] z6655_assgn66558;
    reg [31:0] z2571_assgn2571;
    wire [31:0] i3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6659_assgn6659;
    reg [31:0] z6659_assgn66590;
    reg [31:0] z6659_assgn66591;
    reg [31:0] z6659_assgn66592;
    reg [31:0] z6659_assgn66593;
    reg [31:0] z6659_assgn66594;
    reg [31:0] z6659_assgn66595;
    reg [31:0] z6659_assgn66596;
    reg [31:0] z6659_assgn66597;
    reg [31:0] z6659_assgn66598;
    reg [31:0] z2574_assgn2574;
    reg [31:0] i2_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6663_assgn6663;
    reg [31:0] z6663_assgn66630;
    reg [31:0] z6663_assgn66631;
    reg [31:0] z6663_assgn66632;
    reg [31:0] z6663_assgn66633;
    reg [31:0] z6663_assgn66634;
    reg [31:0] z6663_assgn66635;
    reg [31:0] z6663_assgn66636;
    reg [31:0] z6663_assgn66637;
    reg [31:0] z6663_assgn66638;
    reg [31:0] z2576_assgn2576;
    reg [31:0] i3_comar1_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r00_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m0_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] m2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6701_assgn6701;
    reg [31:0] z6701_assgn67010;
    reg [31:0] z6701_assgn67011;
    reg [31:0] z6701_assgn67012;
    reg [31:0] z6701_assgn67013;
    reg [31:0] z6701_assgn67014;
    reg [31:0] z6701_assgn67015;
    reg [31:0] z6701_assgn67016;
    reg [31:0] z6701_assgn67017;
    reg [31:0] z2611_assgn2611;
    wire [31:0] m3_comar2_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m0_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6707_assgn6707;
    reg [31:0] z6707_assgn67070;
    reg [31:0] z6707_assgn67071;
    reg [31:0] z6707_assgn67072;
    reg [31:0] z6707_assgn67073;
    reg [31:0] z6707_assgn67074;
    reg [31:0] z6707_assgn67075;
    reg [31:0] z6707_assgn67076;
    reg [31:0] z6707_assgn67077;
    reg [31:0] z6707_assgn67078;
    reg [31:0] z2615_assgn2615;
    reg [31:0] m3_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] m2_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6713_assgn6713;
    reg [31:0] z6713_assgn67130;
    reg [31:0] z6713_assgn67131;
    reg [31:0] z6713_assgn67132;
    reg [31:0] z6713_assgn67133;
    reg [31:0] z6713_assgn67134;
    reg [31:0] z6713_assgn67135;
    reg [31:0] z6713_assgn67136;
    reg [31:0] z6713_assgn67137;
    reg [31:0] z6713_assgn67138;
    reg [31:0] z2619_assgn2619;
    wire [31:0] p4_comar2_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6721_assgn6721;
    reg [31:0] z6721_assgn67210;
    reg [31:0] z6721_assgn67211;
    reg [31:0] z6721_assgn67212;
    reg [31:0] z6721_assgn67213;
    reg [31:0] z6721_assgn67214;
    reg [31:0] z6721_assgn67215;
    reg [31:0] z6721_assgn67216;
    reg [31:0] z6721_assgn67217;
    reg [31:0] z6721_assgn67218;
    reg [31:0] z2625_assgn2625;
    wire [31:0] i2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6725_assgn6725;
    reg [31:0] z6725_assgn67250;
    reg [31:0] z6725_assgn67251;
    reg [31:0] z6725_assgn67252;
    reg [31:0] z6725_assgn67253;
    reg [31:0] z6725_assgn67254;
    reg [31:0] z6725_assgn67255;
    reg [31:0] z6725_assgn67256;
    reg [31:0] z6725_assgn67257;
    reg [31:0] z6725_assgn67258;
    reg [31:0] z2627_assgn2627;
    wire [31:0] i3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6729_assgn6729;
    reg [31:0] z6729_assgn67290;
    reg [31:0] z6729_assgn67291;
    reg [31:0] z6729_assgn67292;
    reg [31:0] z6729_assgn67293;
    reg [31:0] z6729_assgn67294;
    reg [31:0] z6729_assgn67295;
    reg [31:0] z6729_assgn67296;
    reg [31:0] z6729_assgn67297;
    reg [31:0] z6729_assgn67298;
    reg [31:0] z2630_assgn2630;
    reg [31:0] i2_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6733_assgn6733;
    reg [31:0] z6733_assgn67330;
    reg [31:0] z6733_assgn67331;
    reg [31:0] z6733_assgn67332;
    reg [31:0] z6733_assgn67333;
    reg [31:0] z6733_assgn67334;
    reg [31:0] z6733_assgn67335;
    reg [31:0] z6733_assgn67336;
    reg [31:0] z6733_assgn67337;
    reg [31:0] z6733_assgn67338;
    reg [31:0] z2632_assgn2632;
    reg [31:0] i3_comar2_G4_mul2_G16_mul1_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0;
    reg [31:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] z6755_assgn6755;
    reg [31:0] z6755_assgn67550;
    reg [31:0] z6755_assgn67551;
    reg [31:0] z6755_assgn67552;
    reg [31:0] z6755_assgn67553;
    reg [31:0] z6755_assgn67554;
    reg [31:0] z6755_assgn67555;
    reg [31:0] z6755_assgn67556;
    reg [31:0] z6755_assgn67557;
    reg [31:0] z6755_assgn67558;
    reg [31:0] z6755_assgn67559;
    reg [31:0] z6755_assgn675510;
    reg [31:0] z2651_assgn2651;
    wire [31:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [31:0] q0_0_G16_mul1_G256_inv0;
    wire [31:0] q1_0_G16_mul1_G256_inv0;
    wire [31:0] q0_G16_mul1_G256_inv0;
    wire [31:0] q1_G16_mul1_G256_inv0;
    wire [31:0] p0ls2_G16_mul1_G256_inv0;
    wire [31:0] z6769_assgn6769;
    reg [31:0] z6769_assgn67690;
    reg [31:0] z6769_assgn67691;
    reg [31:0] z6769_assgn67692;
    reg [31:0] z6769_assgn67693;
    reg [31:0] z6769_assgn67694;
    reg [31:0] z6769_assgn67695;
    reg [31:0] z6769_assgn67696;
    reg [31:0] z6769_assgn67697;
    reg [31:0] z6769_assgn67698;
    reg [31:0] z6769_assgn67699;
    reg [31:0] z6769_assgn676910;
    reg [31:0] z2663_assgn2663;
    wire [31:0] p1ls2_G16_mul1_G256_inv0;
    wire [31:0] p0_G256_inv0;
    wire [31:0] p1_G256_inv0;
    wire [31:0] r00_G16_mul2_G256_inv0;
    wire [31:0] r10_G16_mul2_G256_inv0;
    wire [31:0] r20_G16_mul2_G256_inv0;
    wire [31:0] r30_G16_mul2_G256_inv0;
    wire [31:0] r40_G16_mul2_G256_inv0;
    wire [31:0] r50_G16_mul2_G256_inv0;
    wire [31:0] a0_0_G16_mul2_G256_inv0;
    wire [31:0] z6791_assgn6791;
    reg [31:0] z6791_assgn67910;
    reg [31:0] z6791_assgn67911;
    reg [31:0] z6791_assgn67912;
    reg [31:0] z6791_assgn67913;
    reg [31:0] z6791_assgn67914;
    reg [31:0] z6791_assgn67915;
    reg [31:0] z6791_assgn67916;
    reg [31:0] z6791_assgn67917;
    reg [31:0] z2683_assgn2683;
    wire [31:0] a1_0_G16_mul2_G256_inv0;
    wire [31:0] a0_G16_mul2_G256_inv0;
    wire [31:0] z6797_assgn6797;
    reg [31:0] z6797_assgn67970;
    reg [31:0] z6797_assgn67971;
    reg [31:0] z6797_assgn67972;
    reg [31:0] z6797_assgn67973;
    reg [31:0] z6797_assgn67974;
    reg [31:0] z6797_assgn67975;
    reg [31:0] z6797_assgn67976;
    reg [31:0] z6797_assgn67977;
    reg [31:0] z2687_assgn2687;
    wire [31:0] a1_G16_mul2_G256_inv0;
    wire [31:0] b0_G16_mul2_G256_inv0;
    wire [31:0] z6803_assgn6803;
    reg [31:0] z6803_assgn68030;
    reg [31:0] z6803_assgn68031;
    reg [31:0] z6803_assgn68032;
    reg [31:0] z6803_assgn68033;
    reg [31:0] z6803_assgn68034;
    reg [31:0] z6803_assgn68035;
    reg [31:0] z6803_assgn68036;
    reg [31:0] z6803_assgn68037;
    reg [31:0] z2691_assgn2691;
    wire [31:0] b1_G16_mul2_G256_inv0;
    wire [31:0] c0_0_G16_mul2_G256_inv0;
    wire [31:0] c1_0_G16_mul2_G256_inv0;
    wire [31:0] c0_G16_mul2_G256_inv0;
    wire [31:0] c1_G16_mul2_G256_inv0;
    wire [31:0] d0_G16_mul2_G256_inv0;
    wire [31:0] d1_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G16_mul2_G256_inv0;
    wire [31:0] cxord_0_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G16_mul2_G256_inv0;
    wire [31:0] cxord_1_G16_mul2_G256_inv0;
    wire [31:0] r00_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r10_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r20_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r30_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r40_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r50_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6841_assgn6841;
    reg [31:0] z6841_assgn68410;
    reg [31:0] z6841_assgn68411;
    reg [31:0] z6841_assgn68412;
    reg [31:0] z6841_assgn68413;
    reg [31:0] z6841_assgn68414;
    reg [31:0] z6841_assgn68415;
    reg [31:0] z6841_assgn68416;
    reg [31:0] z6841_assgn68417;
    reg [31:0] z2727_assgn2727;
    wire [31:0] a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6847_assgn6847;
    reg [31:0] z6847_assgn68470;
    reg [31:0] z6847_assgn68471;
    reg [31:0] z6847_assgn68472;
    reg [31:0] z6847_assgn68473;
    reg [31:0] z6847_assgn68474;
    reg [31:0] z6847_assgn68475;
    reg [31:0] z6847_assgn68476;
    reg [31:0] z6847_assgn68477;
    reg [31:0] z2731_assgn2731;
    wire [31:0] a1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6853_assgn6853;
    reg [31:0] z6853_assgn68530;
    reg [31:0] z6853_assgn68531;
    reg [31:0] z6853_assgn68532;
    reg [31:0] z6853_assgn68533;
    reg [31:0] z6853_assgn68534;
    reg [31:0] z6853_assgn68535;
    reg [31:0] z6853_assgn68536;
    reg [31:0] z6853_assgn68537;
    reg [31:0] z2735_assgn2735;
    wire [31:0] b1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] c1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] d1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r00_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m0_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6895_assgn6895;
    reg [31:0] z6895_assgn68950;
    reg [31:0] z6895_assgn68951;
    reg [31:0] z6895_assgn68952;
    reg [31:0] z6895_assgn68953;
    reg [31:0] z6895_assgn68954;
    reg [31:0] z6895_assgn68955;
    reg [31:0] z6895_assgn68956;
    reg [31:0] z6895_assgn68957;
    reg [31:0] z2775_assgn2775;
    wire [31:0] m3_comar0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m0_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6901_assgn6901;
    reg [31:0] z6901_assgn69010;
    reg [31:0] z6901_assgn69011;
    reg [31:0] z6901_assgn69012;
    reg [31:0] z6901_assgn69013;
    reg [31:0] z6901_assgn69014;
    reg [31:0] z6901_assgn69015;
    reg [31:0] z6901_assgn69016;
    reg [31:0] z6901_assgn69017;
    reg [31:0] z6901_assgn69018;
    reg [31:0] z2779_assgn2779;
    reg [31:0] m3_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m2_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6907_assgn6907;
    reg [31:0] z6907_assgn69070;
    reg [31:0] z6907_assgn69071;
    reg [31:0] z6907_assgn69072;
    reg [31:0] z6907_assgn69073;
    reg [31:0] z6907_assgn69074;
    reg [31:0] z6907_assgn69075;
    reg [31:0] z6907_assgn69076;
    reg [31:0] z6907_assgn69077;
    reg [31:0] z6907_assgn69078;
    reg [31:0] z2783_assgn2783;
    wire [31:0] p4_comar0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6915_assgn6915;
    reg [31:0] z6915_assgn69150;
    reg [31:0] z6915_assgn69151;
    reg [31:0] z6915_assgn69152;
    reg [31:0] z6915_assgn69153;
    reg [31:0] z6915_assgn69154;
    reg [31:0] z6915_assgn69155;
    reg [31:0] z6915_assgn69156;
    reg [31:0] z6915_assgn69157;
    reg [31:0] z6915_assgn69158;
    reg [31:0] z2789_assgn2789;
    wire [31:0] i2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6919_assgn6919;
    reg [31:0] z6919_assgn69190;
    reg [31:0] z6919_assgn69191;
    reg [31:0] z6919_assgn69192;
    reg [31:0] z6919_assgn69193;
    reg [31:0] z6919_assgn69194;
    reg [31:0] z6919_assgn69195;
    reg [31:0] z6919_assgn69196;
    reg [31:0] z6919_assgn69197;
    reg [31:0] z6919_assgn69198;
    reg [31:0] z2791_assgn2791;
    wire [31:0] i3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6923_assgn6923;
    reg [31:0] z6923_assgn69230;
    reg [31:0] z6923_assgn69231;
    reg [31:0] z6923_assgn69232;
    reg [31:0] z6923_assgn69233;
    reg [31:0] z6923_assgn69234;
    reg [31:0] z6923_assgn69235;
    reg [31:0] z6923_assgn69236;
    reg [31:0] z6923_assgn69237;
    reg [31:0] z6923_assgn69238;
    reg [31:0] z2794_assgn2794;
    reg [31:0] i2_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6927_assgn6927;
    reg [31:0] z6927_assgn69270;
    reg [31:0] z6927_assgn69271;
    reg [31:0] z6927_assgn69272;
    reg [31:0] z6927_assgn69273;
    reg [31:0] z6927_assgn69274;
    reg [31:0] z6927_assgn69275;
    reg [31:0] z6927_assgn69276;
    reg [31:0] z6927_assgn69277;
    reg [31:0] z6927_assgn69278;
    reg [31:0] z2796_assgn2796;
    reg [31:0] i3_comar0_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] e0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] e1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r00_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m0_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6961_assgn6961;
    reg [31:0] z6961_assgn69610;
    reg [31:0] z6961_assgn69611;
    reg [31:0] z6961_assgn69612;
    reg [31:0] z6961_assgn69613;
    reg [31:0] z6961_assgn69614;
    reg [31:0] z6961_assgn69615;
    reg [31:0] z6961_assgn69616;
    reg [31:0] z6961_assgn69617;
    reg [31:0] z2827_assgn2827;
    wire [31:0] m3_comar1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m0_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6967_assgn6967;
    reg [31:0] z6967_assgn69670;
    reg [31:0] z6967_assgn69671;
    reg [31:0] z6967_assgn69672;
    reg [31:0] z6967_assgn69673;
    reg [31:0] z6967_assgn69674;
    reg [31:0] z6967_assgn69675;
    reg [31:0] z6967_assgn69676;
    reg [31:0] z6967_assgn69677;
    reg [31:0] z6967_assgn69678;
    reg [31:0] z2831_assgn2831;
    reg [31:0] m3_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m2_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6973_assgn6973;
    reg [31:0] z6973_assgn69730;
    reg [31:0] z6973_assgn69731;
    reg [31:0] z6973_assgn69732;
    reg [31:0] z6973_assgn69733;
    reg [31:0] z6973_assgn69734;
    reg [31:0] z6973_assgn69735;
    reg [31:0] z6973_assgn69736;
    reg [31:0] z6973_assgn69737;
    reg [31:0] z6973_assgn69738;
    reg [31:0] z2835_assgn2835;
    wire [31:0] p4_comar1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6981_assgn6981;
    reg [31:0] z6981_assgn69810;
    reg [31:0] z6981_assgn69811;
    reg [31:0] z6981_assgn69812;
    reg [31:0] z6981_assgn69813;
    reg [31:0] z6981_assgn69814;
    reg [31:0] z6981_assgn69815;
    reg [31:0] z6981_assgn69816;
    reg [31:0] z6981_assgn69817;
    reg [31:0] z6981_assgn69818;
    reg [31:0] z2841_assgn2841;
    wire [31:0] i2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6985_assgn6985;
    reg [31:0] z6985_assgn69850;
    reg [31:0] z6985_assgn69851;
    reg [31:0] z6985_assgn69852;
    reg [31:0] z6985_assgn69853;
    reg [31:0] z6985_assgn69854;
    reg [31:0] z6985_assgn69855;
    reg [31:0] z6985_assgn69856;
    reg [31:0] z6985_assgn69857;
    reg [31:0] z6985_assgn69858;
    reg [31:0] z2843_assgn2843;
    wire [31:0] i3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6989_assgn6989;
    reg [31:0] z6989_assgn69890;
    reg [31:0] z6989_assgn69891;
    reg [31:0] z6989_assgn69892;
    reg [31:0] z6989_assgn69893;
    reg [31:0] z6989_assgn69894;
    reg [31:0] z6989_assgn69895;
    reg [31:0] z6989_assgn69896;
    reg [31:0] z6989_assgn69897;
    reg [31:0] z6989_assgn69898;
    reg [31:0] z2846_assgn2846;
    reg [31:0] i2_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z6993_assgn6993;
    reg [31:0] z6993_assgn69930;
    reg [31:0] z6993_assgn69931;
    reg [31:0] z6993_assgn69932;
    reg [31:0] z6993_assgn69933;
    reg [31:0] z6993_assgn69934;
    reg [31:0] z6993_assgn69935;
    reg [31:0] z6993_assgn69936;
    reg [31:0] z6993_assgn69937;
    reg [31:0] z6993_assgn69938;
    reg [31:0] z2848_assgn2848;
    reg [31:0] i3_comar1_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r00_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m0_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] m2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7031_assgn7031;
    reg [31:0] z7031_assgn70310;
    reg [31:0] z7031_assgn70311;
    reg [31:0] z7031_assgn70312;
    reg [31:0] z7031_assgn70313;
    reg [31:0] z7031_assgn70314;
    reg [31:0] z7031_assgn70315;
    reg [31:0] z7031_assgn70316;
    reg [31:0] z7031_assgn70317;
    reg [31:0] z2883_assgn2883;
    wire [31:0] m3_comar2_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m0_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7037_assgn7037;
    reg [31:0] z7037_assgn70370;
    reg [31:0] z7037_assgn70371;
    reg [31:0] z7037_assgn70372;
    reg [31:0] z7037_assgn70373;
    reg [31:0] z7037_assgn70374;
    reg [31:0] z7037_assgn70375;
    reg [31:0] z7037_assgn70376;
    reg [31:0] z7037_assgn70377;
    reg [31:0] z7037_assgn70378;
    reg [31:0] z2887_assgn2887;
    reg [31:0] m3_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] m2_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7043_assgn7043;
    reg [31:0] z7043_assgn70430;
    reg [31:0] z7043_assgn70431;
    reg [31:0] z7043_assgn70432;
    reg [31:0] z7043_assgn70433;
    reg [31:0] z7043_assgn70434;
    reg [31:0] z7043_assgn70435;
    reg [31:0] z7043_assgn70436;
    reg [31:0] z7043_assgn70437;
    reg [31:0] z7043_assgn70438;
    reg [31:0] z2891_assgn2891;
    wire [31:0] p4_comar2_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7051_assgn7051;
    reg [31:0] z7051_assgn70510;
    reg [31:0] z7051_assgn70511;
    reg [31:0] z7051_assgn70512;
    reg [31:0] z7051_assgn70513;
    reg [31:0] z7051_assgn70514;
    reg [31:0] z7051_assgn70515;
    reg [31:0] z7051_assgn70516;
    reg [31:0] z7051_assgn70517;
    reg [31:0] z7051_assgn70518;
    reg [31:0] z2897_assgn2897;
    wire [31:0] i2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7055_assgn7055;
    reg [31:0] z7055_assgn70550;
    reg [31:0] z7055_assgn70551;
    reg [31:0] z7055_assgn70552;
    reg [31:0] z7055_assgn70553;
    reg [31:0] z7055_assgn70554;
    reg [31:0] z7055_assgn70555;
    reg [31:0] z7055_assgn70556;
    reg [31:0] z7055_assgn70557;
    reg [31:0] z7055_assgn70558;
    reg [31:0] z2899_assgn2899;
    wire [31:0] i3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7059_assgn7059;
    reg [31:0] z7059_assgn70590;
    reg [31:0] z7059_assgn70591;
    reg [31:0] z7059_assgn70592;
    reg [31:0] z7059_assgn70593;
    reg [31:0] z7059_assgn70594;
    reg [31:0] z7059_assgn70595;
    reg [31:0] z7059_assgn70596;
    reg [31:0] z7059_assgn70597;
    reg [31:0] z7059_assgn70598;
    reg [31:0] z2902_assgn2902;
    reg [31:0] i2_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7063_assgn7063;
    reg [31:0] z7063_assgn70630;
    reg [31:0] z7063_assgn70631;
    reg [31:0] z7063_assgn70632;
    reg [31:0] z7063_assgn70633;
    reg [31:0] z7063_assgn70634;
    reg [31:0] z7063_assgn70635;
    reg [31:0] z7063_assgn70636;
    reg [31:0] z7063_assgn70637;
    reg [31:0] z7063_assgn70638;
    reg [31:0] z2904_assgn2904;
    reg [31:0] i3_comar2_G4_mul0_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0;
    reg [31:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] z7085_assgn7085;
    reg [31:0] z7085_assgn70850;
    reg [31:0] z7085_assgn70851;
    reg [31:0] z7085_assgn70852;
    reg [31:0] z7085_assgn70853;
    reg [31:0] z7085_assgn70854;
    reg [31:0] z7085_assgn70855;
    reg [31:0] z7085_assgn70856;
    reg [31:0] z7085_assgn70857;
    reg [31:0] z7085_assgn70858;
    reg [31:0] z7085_assgn70859;
    reg [31:0] z7085_assgn708510;
    reg [31:0] z2923_assgn2923;
    wire [31:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [31:0] e0_G16_mul2_G256_inv0;
    wire [31:0] e1_G16_mul2_G256_inv0;
    wire [31:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z7095_assgn7095;
    reg [31:0] z7095_assgn70950;
    reg [31:0] z7095_assgn70951;
    reg [31:0] z7095_assgn70952;
    reg [31:0] z7095_assgn70953;
    reg [31:0] z7095_assgn70954;
    reg [31:0] z7095_assgn70955;
    reg [31:0] z7095_assgn70956;
    reg [31:0] z7095_assgn70957;
    reg [31:0] z7095_assgn70958;
    reg [31:0] z7095_assgn70959;
    reg [31:0] z7095_assgn709510;
    reg [31:0] z2931_assgn2931;
    wire [31:0] a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z7101_assgn7101;
    reg [31:0] z7101_assgn71010;
    reg [31:0] z7101_assgn71011;
    reg [31:0] z7101_assgn71012;
    reg [31:0] z7101_assgn71013;
    reg [31:0] z7101_assgn71014;
    reg [31:0] z7101_assgn71015;
    reg [31:0] z7101_assgn71016;
    reg [31:0] z7101_assgn71017;
    reg [31:0] z7101_assgn71018;
    reg [31:0] z7101_assgn71019;
    reg [31:0] z7101_assgn710110;
    reg [31:0] z2935_assgn2935;
    wire [31:0] a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z7107_assgn7107;
    reg [31:0] z7107_assgn71070;
    reg [31:0] z7107_assgn71071;
    reg [31:0] z7107_assgn71072;
    reg [31:0] z7107_assgn71073;
    reg [31:0] z7107_assgn71074;
    reg [31:0] z7107_assgn71075;
    reg [31:0] z7107_assgn71076;
    reg [31:0] z7107_assgn71077;
    reg [31:0] z7107_assgn71078;
    reg [31:0] z7107_assgn71079;
    reg [31:0] z7107_assgn710710;
    reg [31:0] z2939_assgn2939;
    wire [31:0] b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] z7119_assgn7119;
    reg [31:0] z7119_assgn71190;
    reg [31:0] z7119_assgn71191;
    reg [31:0] z7119_assgn71192;
    reg [31:0] z7119_assgn71193;
    reg [31:0] z7119_assgn71194;
    reg [31:0] z7119_assgn71195;
    reg [31:0] z7119_assgn71196;
    reg [31:0] z7119_assgn71197;
    reg [31:0] z7119_assgn71198;
    reg [31:0] z7119_assgn71199;
    reg [31:0] z7119_assgn711910;
    reg [31:0] z2949_assgn2949;
    wire [31:0] p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [31:0] e01_G16_mul2_G256_inv0;
    wire [31:0] e11_G16_mul2_G256_inv0;
    wire [31:0] r00_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r10_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r20_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r30_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r40_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r50_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7143_assgn7143;
    reg [31:0] z7143_assgn71430;
    reg [31:0] z7143_assgn71431;
    reg [31:0] z7143_assgn71432;
    reg [31:0] z7143_assgn71433;
    reg [31:0] z7143_assgn71434;
    reg [31:0] z7143_assgn71435;
    reg [31:0] z7143_assgn71436;
    reg [31:0] z7143_assgn71437;
    reg [31:0] z2971_assgn2971;
    wire [31:0] a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7149_assgn7149;
    reg [31:0] z7149_assgn71490;
    reg [31:0] z7149_assgn71491;
    reg [31:0] z7149_assgn71492;
    reg [31:0] z7149_assgn71493;
    reg [31:0] z7149_assgn71494;
    reg [31:0] z7149_assgn71495;
    reg [31:0] z7149_assgn71496;
    reg [31:0] z7149_assgn71497;
    reg [31:0] z2975_assgn2975;
    wire [31:0] a1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7155_assgn7155;
    reg [31:0] z7155_assgn71550;
    reg [31:0] z7155_assgn71551;
    reg [31:0] z7155_assgn71552;
    reg [31:0] z7155_assgn71553;
    reg [31:0] z7155_assgn71554;
    reg [31:0] z7155_assgn71555;
    reg [31:0] z7155_assgn71556;
    reg [31:0] z7155_assgn71557;
    reg [31:0] z2979_assgn2979;
    wire [31:0] b1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] c1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] d1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r00_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m0_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7197_assgn7197;
    reg [31:0] z7197_assgn71970;
    reg [31:0] z7197_assgn71971;
    reg [31:0] z7197_assgn71972;
    reg [31:0] z7197_assgn71973;
    reg [31:0] z7197_assgn71974;
    reg [31:0] z7197_assgn71975;
    reg [31:0] z7197_assgn71976;
    reg [31:0] z7197_assgn71977;
    reg [31:0] z3019_assgn3019;
    wire [31:0] m3_comar0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m0_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7203_assgn7203;
    reg [31:0] z7203_assgn72030;
    reg [31:0] z7203_assgn72031;
    reg [31:0] z7203_assgn72032;
    reg [31:0] z7203_assgn72033;
    reg [31:0] z7203_assgn72034;
    reg [31:0] z7203_assgn72035;
    reg [31:0] z7203_assgn72036;
    reg [31:0] z7203_assgn72037;
    reg [31:0] z7203_assgn72038;
    reg [31:0] z3023_assgn3023;
    reg [31:0] m3_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m2_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7209_assgn7209;
    reg [31:0] z7209_assgn72090;
    reg [31:0] z7209_assgn72091;
    reg [31:0] z7209_assgn72092;
    reg [31:0] z7209_assgn72093;
    reg [31:0] z7209_assgn72094;
    reg [31:0] z7209_assgn72095;
    reg [31:0] z7209_assgn72096;
    reg [31:0] z7209_assgn72097;
    reg [31:0] z7209_assgn72098;
    reg [31:0] z3027_assgn3027;
    wire [31:0] p4_comar0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7217_assgn7217;
    reg [31:0] z7217_assgn72170;
    reg [31:0] z7217_assgn72171;
    reg [31:0] z7217_assgn72172;
    reg [31:0] z7217_assgn72173;
    reg [31:0] z7217_assgn72174;
    reg [31:0] z7217_assgn72175;
    reg [31:0] z7217_assgn72176;
    reg [31:0] z7217_assgn72177;
    reg [31:0] z7217_assgn72178;
    reg [31:0] z3033_assgn3033;
    wire [31:0] i2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7221_assgn7221;
    reg [31:0] z7221_assgn72210;
    reg [31:0] z7221_assgn72211;
    reg [31:0] z7221_assgn72212;
    reg [31:0] z7221_assgn72213;
    reg [31:0] z7221_assgn72214;
    reg [31:0] z7221_assgn72215;
    reg [31:0] z7221_assgn72216;
    reg [31:0] z7221_assgn72217;
    reg [31:0] z7221_assgn72218;
    reg [31:0] z3035_assgn3035;
    wire [31:0] i3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7225_assgn7225;
    reg [31:0] z7225_assgn72250;
    reg [31:0] z7225_assgn72251;
    reg [31:0] z7225_assgn72252;
    reg [31:0] z7225_assgn72253;
    reg [31:0] z7225_assgn72254;
    reg [31:0] z7225_assgn72255;
    reg [31:0] z7225_assgn72256;
    reg [31:0] z7225_assgn72257;
    reg [31:0] z7225_assgn72258;
    reg [31:0] z3038_assgn3038;
    reg [31:0] i2_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7229_assgn7229;
    reg [31:0] z7229_assgn72290;
    reg [31:0] z7229_assgn72291;
    reg [31:0] z7229_assgn72292;
    reg [31:0] z7229_assgn72293;
    reg [31:0] z7229_assgn72294;
    reg [31:0] z7229_assgn72295;
    reg [31:0] z7229_assgn72296;
    reg [31:0] z7229_assgn72297;
    reg [31:0] z7229_assgn72298;
    reg [31:0] z3040_assgn3040;
    reg [31:0] i3_comar0_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] e0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] e1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r00_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m0_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7263_assgn7263;
    reg [31:0] z7263_assgn72630;
    reg [31:0] z7263_assgn72631;
    reg [31:0] z7263_assgn72632;
    reg [31:0] z7263_assgn72633;
    reg [31:0] z7263_assgn72634;
    reg [31:0] z7263_assgn72635;
    reg [31:0] z7263_assgn72636;
    reg [31:0] z7263_assgn72637;
    reg [31:0] z3071_assgn3071;
    wire [31:0] m3_comar1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m0_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7269_assgn7269;
    reg [31:0] z7269_assgn72690;
    reg [31:0] z7269_assgn72691;
    reg [31:0] z7269_assgn72692;
    reg [31:0] z7269_assgn72693;
    reg [31:0] z7269_assgn72694;
    reg [31:0] z7269_assgn72695;
    reg [31:0] z7269_assgn72696;
    reg [31:0] z7269_assgn72697;
    reg [31:0] z7269_assgn72698;
    reg [31:0] z3075_assgn3075;
    reg [31:0] m3_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m2_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7275_assgn7275;
    reg [31:0] z7275_assgn72750;
    reg [31:0] z7275_assgn72751;
    reg [31:0] z7275_assgn72752;
    reg [31:0] z7275_assgn72753;
    reg [31:0] z7275_assgn72754;
    reg [31:0] z7275_assgn72755;
    reg [31:0] z7275_assgn72756;
    reg [31:0] z7275_assgn72757;
    reg [31:0] z7275_assgn72758;
    reg [31:0] z3079_assgn3079;
    wire [31:0] p4_comar1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7283_assgn7283;
    reg [31:0] z7283_assgn72830;
    reg [31:0] z7283_assgn72831;
    reg [31:0] z7283_assgn72832;
    reg [31:0] z7283_assgn72833;
    reg [31:0] z7283_assgn72834;
    reg [31:0] z7283_assgn72835;
    reg [31:0] z7283_assgn72836;
    reg [31:0] z7283_assgn72837;
    reg [31:0] z7283_assgn72838;
    reg [31:0] z3085_assgn3085;
    wire [31:0] i2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7287_assgn7287;
    reg [31:0] z7287_assgn72870;
    reg [31:0] z7287_assgn72871;
    reg [31:0] z7287_assgn72872;
    reg [31:0] z7287_assgn72873;
    reg [31:0] z7287_assgn72874;
    reg [31:0] z7287_assgn72875;
    reg [31:0] z7287_assgn72876;
    reg [31:0] z7287_assgn72877;
    reg [31:0] z7287_assgn72878;
    reg [31:0] z3087_assgn3087;
    wire [31:0] i3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7291_assgn7291;
    reg [31:0] z7291_assgn72910;
    reg [31:0] z7291_assgn72911;
    reg [31:0] z7291_assgn72912;
    reg [31:0] z7291_assgn72913;
    reg [31:0] z7291_assgn72914;
    reg [31:0] z7291_assgn72915;
    reg [31:0] z7291_assgn72916;
    reg [31:0] z7291_assgn72917;
    reg [31:0] z7291_assgn72918;
    reg [31:0] z3090_assgn3090;
    reg [31:0] i2_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7295_assgn7295;
    reg [31:0] z7295_assgn72950;
    reg [31:0] z7295_assgn72951;
    reg [31:0] z7295_assgn72952;
    reg [31:0] z7295_assgn72953;
    reg [31:0] z7295_assgn72954;
    reg [31:0] z7295_assgn72955;
    reg [31:0] z7295_assgn72956;
    reg [31:0] z7295_assgn72957;
    reg [31:0] z7295_assgn72958;
    reg [31:0] z3092_assgn3092;
    reg [31:0] i3_comar1_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r00_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m0_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] m2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7333_assgn7333;
    reg [31:0] z7333_assgn73330;
    reg [31:0] z7333_assgn73331;
    reg [31:0] z7333_assgn73332;
    reg [31:0] z7333_assgn73333;
    reg [31:0] z7333_assgn73334;
    reg [31:0] z7333_assgn73335;
    reg [31:0] z7333_assgn73336;
    reg [31:0] z7333_assgn73337;
    reg [31:0] z3127_assgn3127;
    wire [31:0] m3_comar2_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m0_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7339_assgn7339;
    reg [31:0] z7339_assgn73390;
    reg [31:0] z7339_assgn73391;
    reg [31:0] z7339_assgn73392;
    reg [31:0] z7339_assgn73393;
    reg [31:0] z7339_assgn73394;
    reg [31:0] z7339_assgn73395;
    reg [31:0] z7339_assgn73396;
    reg [31:0] z7339_assgn73397;
    reg [31:0] z7339_assgn73398;
    reg [31:0] z3131_assgn3131;
    reg [31:0] m3_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] m2_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7345_assgn7345;
    reg [31:0] z7345_assgn73450;
    reg [31:0] z7345_assgn73451;
    reg [31:0] z7345_assgn73452;
    reg [31:0] z7345_assgn73453;
    reg [31:0] z7345_assgn73454;
    reg [31:0] z7345_assgn73455;
    reg [31:0] z7345_assgn73456;
    reg [31:0] z7345_assgn73457;
    reg [31:0] z7345_assgn73458;
    reg [31:0] z3135_assgn3135;
    wire [31:0] p4_comar2_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7353_assgn7353;
    reg [31:0] z7353_assgn73530;
    reg [31:0] z7353_assgn73531;
    reg [31:0] z7353_assgn73532;
    reg [31:0] z7353_assgn73533;
    reg [31:0] z7353_assgn73534;
    reg [31:0] z7353_assgn73535;
    reg [31:0] z7353_assgn73536;
    reg [31:0] z7353_assgn73537;
    reg [31:0] z7353_assgn73538;
    reg [31:0] z3141_assgn3141;
    wire [31:0] i2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7357_assgn7357;
    reg [31:0] z7357_assgn73570;
    reg [31:0] z7357_assgn73571;
    reg [31:0] z7357_assgn73572;
    reg [31:0] z7357_assgn73573;
    reg [31:0] z7357_assgn73574;
    reg [31:0] z7357_assgn73575;
    reg [31:0] z7357_assgn73576;
    reg [31:0] z7357_assgn73577;
    reg [31:0] z7357_assgn73578;
    reg [31:0] z3143_assgn3143;
    wire [31:0] i3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7361_assgn7361;
    reg [31:0] z7361_assgn73610;
    reg [31:0] z7361_assgn73611;
    reg [31:0] z7361_assgn73612;
    reg [31:0] z7361_assgn73613;
    reg [31:0] z7361_assgn73614;
    reg [31:0] z7361_assgn73615;
    reg [31:0] z7361_assgn73616;
    reg [31:0] z7361_assgn73617;
    reg [31:0] z7361_assgn73618;
    reg [31:0] z3146_assgn3146;
    reg [31:0] i2_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7365_assgn7365;
    reg [31:0] z7365_assgn73650;
    reg [31:0] z7365_assgn73651;
    reg [31:0] z7365_assgn73652;
    reg [31:0] z7365_assgn73653;
    reg [31:0] z7365_assgn73654;
    reg [31:0] z7365_assgn73655;
    reg [31:0] z7365_assgn73656;
    reg [31:0] z7365_assgn73657;
    reg [31:0] z7365_assgn73658;
    reg [31:0] z3148_assgn3148;
    reg [31:0] i3_comar2_G4_mul1_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0;
    reg [31:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] z7387_assgn7387;
    reg [31:0] z7387_assgn73870;
    reg [31:0] z7387_assgn73871;
    reg [31:0] z7387_assgn73872;
    reg [31:0] z7387_assgn73873;
    reg [31:0] z7387_assgn73874;
    reg [31:0] z7387_assgn73875;
    reg [31:0] z7387_assgn73876;
    reg [31:0] z7387_assgn73877;
    reg [31:0] z7387_assgn73878;
    reg [31:0] z7387_assgn73879;
    reg [31:0] z7387_assgn738710;
    reg [31:0] z3167_assgn3167;
    wire [31:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [31:0] p0_0_G16_mul2_G256_inv0;
    wire [31:0] p1_0_G16_mul2_G256_inv0;
    wire [31:0] p0_G16_mul2_G256_inv0;
    wire [31:0] p1_G16_mul2_G256_inv0;
    wire [31:0] r00_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r10_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r20_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r30_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r40_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r50_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7413_assgn7413;
    reg [31:0] z7413_assgn74130;
    reg [31:0] z7413_assgn74131;
    reg [31:0] z7413_assgn74132;
    reg [31:0] z7413_assgn74133;
    reg [31:0] z7413_assgn74134;
    reg [31:0] z7413_assgn74135;
    reg [31:0] z7413_assgn74136;
    reg [31:0] z7413_assgn74137;
    reg [31:0] z3191_assgn3191;
    wire [31:0] a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7419_assgn7419;
    reg [31:0] z7419_assgn74190;
    reg [31:0] z7419_assgn74191;
    reg [31:0] z7419_assgn74192;
    reg [31:0] z7419_assgn74193;
    reg [31:0] z7419_assgn74194;
    reg [31:0] z7419_assgn74195;
    reg [31:0] z7419_assgn74196;
    reg [31:0] z7419_assgn74197;
    reg [31:0] z3195_assgn3195;
    wire [31:0] a1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7425_assgn7425;
    reg [31:0] z7425_assgn74250;
    reg [31:0] z7425_assgn74251;
    reg [31:0] z7425_assgn74252;
    reg [31:0] z7425_assgn74253;
    reg [31:0] z7425_assgn74254;
    reg [31:0] z7425_assgn74255;
    reg [31:0] z7425_assgn74256;
    reg [31:0] z7425_assgn74257;
    reg [31:0] z3199_assgn3199;
    wire [31:0] b1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] c1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] d1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] axorb_1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r00_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m0_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7467_assgn7467;
    reg [31:0] z7467_assgn74670;
    reg [31:0] z7467_assgn74671;
    reg [31:0] z7467_assgn74672;
    reg [31:0] z7467_assgn74673;
    reg [31:0] z7467_assgn74674;
    reg [31:0] z7467_assgn74675;
    reg [31:0] z7467_assgn74676;
    reg [31:0] z7467_assgn74677;
    reg [31:0] z3239_assgn3239;
    wire [31:0] m3_comar0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m0_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7473_assgn7473;
    reg [31:0] z7473_assgn74730;
    reg [31:0] z7473_assgn74731;
    reg [31:0] z7473_assgn74732;
    reg [31:0] z7473_assgn74733;
    reg [31:0] z7473_assgn74734;
    reg [31:0] z7473_assgn74735;
    reg [31:0] z7473_assgn74736;
    reg [31:0] z7473_assgn74737;
    reg [31:0] z7473_assgn74738;
    reg [31:0] z3243_assgn3243;
    reg [31:0] m3_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m2_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7479_assgn7479;
    reg [31:0] z7479_assgn74790;
    reg [31:0] z7479_assgn74791;
    reg [31:0] z7479_assgn74792;
    reg [31:0] z7479_assgn74793;
    reg [31:0] z7479_assgn74794;
    reg [31:0] z7479_assgn74795;
    reg [31:0] z7479_assgn74796;
    reg [31:0] z7479_assgn74797;
    reg [31:0] z7479_assgn74798;
    reg [31:0] z3247_assgn3247;
    wire [31:0] p4_comar0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7487_assgn7487;
    reg [31:0] z7487_assgn74870;
    reg [31:0] z7487_assgn74871;
    reg [31:0] z7487_assgn74872;
    reg [31:0] z7487_assgn74873;
    reg [31:0] z7487_assgn74874;
    reg [31:0] z7487_assgn74875;
    reg [31:0] z7487_assgn74876;
    reg [31:0] z7487_assgn74877;
    reg [31:0] z7487_assgn74878;
    reg [31:0] z3253_assgn3253;
    wire [31:0] i2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7491_assgn7491;
    reg [31:0] z7491_assgn74910;
    reg [31:0] z7491_assgn74911;
    reg [31:0] z7491_assgn74912;
    reg [31:0] z7491_assgn74913;
    reg [31:0] z7491_assgn74914;
    reg [31:0] z7491_assgn74915;
    reg [31:0] z7491_assgn74916;
    reg [31:0] z7491_assgn74917;
    reg [31:0] z7491_assgn74918;
    reg [31:0] z3255_assgn3255;
    wire [31:0] i3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7495_assgn7495;
    reg [31:0] z7495_assgn74950;
    reg [31:0] z7495_assgn74951;
    reg [31:0] z7495_assgn74952;
    reg [31:0] z7495_assgn74953;
    reg [31:0] z7495_assgn74954;
    reg [31:0] z7495_assgn74955;
    reg [31:0] z7495_assgn74956;
    reg [31:0] z7495_assgn74957;
    reg [31:0] z7495_assgn74958;
    reg [31:0] z3258_assgn3258;
    reg [31:0] i2_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7499_assgn7499;
    reg [31:0] z7499_assgn74990;
    reg [31:0] z7499_assgn74991;
    reg [31:0] z7499_assgn74992;
    reg [31:0] z7499_assgn74993;
    reg [31:0] z7499_assgn74994;
    reg [31:0] z7499_assgn74995;
    reg [31:0] z7499_assgn74996;
    reg [31:0] z7499_assgn74997;
    reg [31:0] z7499_assgn74998;
    reg [31:0] z3260_assgn3260;
    reg [31:0] i3_comar0_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] e0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] e1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r00_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m0_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7533_assgn7533;
    reg [31:0] z7533_assgn75330;
    reg [31:0] z7533_assgn75331;
    reg [31:0] z7533_assgn75332;
    reg [31:0] z7533_assgn75333;
    reg [31:0] z7533_assgn75334;
    reg [31:0] z7533_assgn75335;
    reg [31:0] z7533_assgn75336;
    reg [31:0] z7533_assgn75337;
    reg [31:0] z3291_assgn3291;
    wire [31:0] m3_comar1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m0_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7539_assgn7539;
    reg [31:0] z7539_assgn75390;
    reg [31:0] z7539_assgn75391;
    reg [31:0] z7539_assgn75392;
    reg [31:0] z7539_assgn75393;
    reg [31:0] z7539_assgn75394;
    reg [31:0] z7539_assgn75395;
    reg [31:0] z7539_assgn75396;
    reg [31:0] z7539_assgn75397;
    reg [31:0] z7539_assgn75398;
    reg [31:0] z3295_assgn3295;
    reg [31:0] m3_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m2_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7545_assgn7545;
    reg [31:0] z7545_assgn75450;
    reg [31:0] z7545_assgn75451;
    reg [31:0] z7545_assgn75452;
    reg [31:0] z7545_assgn75453;
    reg [31:0] z7545_assgn75454;
    reg [31:0] z7545_assgn75455;
    reg [31:0] z7545_assgn75456;
    reg [31:0] z7545_assgn75457;
    reg [31:0] z7545_assgn75458;
    reg [31:0] z3299_assgn3299;
    wire [31:0] p4_comar1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7553_assgn7553;
    reg [31:0] z7553_assgn75530;
    reg [31:0] z7553_assgn75531;
    reg [31:0] z7553_assgn75532;
    reg [31:0] z7553_assgn75533;
    reg [31:0] z7553_assgn75534;
    reg [31:0] z7553_assgn75535;
    reg [31:0] z7553_assgn75536;
    reg [31:0] z7553_assgn75537;
    reg [31:0] z7553_assgn75538;
    reg [31:0] z3305_assgn3305;
    wire [31:0] i2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7557_assgn7557;
    reg [31:0] z7557_assgn75570;
    reg [31:0] z7557_assgn75571;
    reg [31:0] z7557_assgn75572;
    reg [31:0] z7557_assgn75573;
    reg [31:0] z7557_assgn75574;
    reg [31:0] z7557_assgn75575;
    reg [31:0] z7557_assgn75576;
    reg [31:0] z7557_assgn75577;
    reg [31:0] z7557_assgn75578;
    reg [31:0] z3307_assgn3307;
    wire [31:0] i3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7561_assgn7561;
    reg [31:0] z7561_assgn75610;
    reg [31:0] z7561_assgn75611;
    reg [31:0] z7561_assgn75612;
    reg [31:0] z7561_assgn75613;
    reg [31:0] z7561_assgn75614;
    reg [31:0] z7561_assgn75615;
    reg [31:0] z7561_assgn75616;
    reg [31:0] z7561_assgn75617;
    reg [31:0] z7561_assgn75618;
    reg [31:0] z3310_assgn3310;
    reg [31:0] i2_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7565_assgn7565;
    reg [31:0] z7565_assgn75650;
    reg [31:0] z7565_assgn75651;
    reg [31:0] z7565_assgn75652;
    reg [31:0] z7565_assgn75653;
    reg [31:0] z7565_assgn75654;
    reg [31:0] z7565_assgn75655;
    reg [31:0] z7565_assgn75656;
    reg [31:0] z7565_assgn75657;
    reg [31:0] z7565_assgn75658;
    reg [31:0] z3312_assgn3312;
    reg [31:0] i3_comar1_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r00_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r0_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r1_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r2_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] r3_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m0_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] m2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7603_assgn7603;
    reg [31:0] z7603_assgn76030;
    reg [31:0] z7603_assgn76031;
    reg [31:0] z7603_assgn76032;
    reg [31:0] z7603_assgn76033;
    reg [31:0] z7603_assgn76034;
    reg [31:0] z7603_assgn76035;
    reg [31:0] z7603_assgn76036;
    reg [31:0] z7603_assgn76037;
    reg [31:0] z3347_assgn3347;
    wire [31:0] m3_comar2_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m0_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    reg [31:0] m1_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7609_assgn7609;
    reg [31:0] z7609_assgn76090;
    reg [31:0] z7609_assgn76091;
    reg [31:0] z7609_assgn76092;
    reg [31:0] z7609_assgn76093;
    reg [31:0] z7609_assgn76094;
    reg [31:0] z7609_assgn76095;
    reg [31:0] z7609_assgn76096;
    reg [31:0] z7609_assgn76097;
    reg [31:0] z7609_assgn76098;
    reg [31:0] z3351_assgn3351;
    reg [31:0] m3_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p3_comar2_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] m2_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] p1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7615_assgn7615;
    reg [31:0] z7615_assgn76150;
    reg [31:0] z7615_assgn76151;
    reg [31:0] z7615_assgn76152;
    reg [31:0] z7615_assgn76153;
    reg [31:0] z7615_assgn76154;
    reg [31:0] z7615_assgn76155;
    reg [31:0] z7615_assgn76156;
    reg [31:0] z7615_assgn76157;
    reg [31:0] z7615_assgn76158;
    reg [31:0] z3355_assgn3355;
    wire [31:0] p4_comar2_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r0_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0_comar2_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] r1_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7623_assgn7623;
    reg [31:0] z7623_assgn76230;
    reg [31:0] z7623_assgn76231;
    reg [31:0] z7623_assgn76232;
    reg [31:0] z7623_assgn76233;
    reg [31:0] z7623_assgn76234;
    reg [31:0] z7623_assgn76235;
    reg [31:0] z7623_assgn76236;
    reg [31:0] z7623_assgn76237;
    reg [31:0] z7623_assgn76238;
    reg [31:0] z3361_assgn3361;
    wire [31:0] i2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7627_assgn7627;
    reg [31:0] z7627_assgn76270;
    reg [31:0] z7627_assgn76271;
    reg [31:0] z7627_assgn76272;
    reg [31:0] z7627_assgn76273;
    reg [31:0] z7627_assgn76274;
    reg [31:0] z7627_assgn76275;
    reg [31:0] z7627_assgn76276;
    reg [31:0] z7627_assgn76277;
    reg [31:0] z7627_assgn76278;
    reg [31:0] z3363_assgn3363;
    wire [31:0] i3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7631_assgn7631;
    reg [31:0] z7631_assgn76310;
    reg [31:0] z7631_assgn76311;
    reg [31:0] z7631_assgn76312;
    reg [31:0] z7631_assgn76313;
    reg [31:0] z7631_assgn76314;
    reg [31:0] z7631_assgn76315;
    reg [31:0] z7631_assgn76316;
    reg [31:0] z7631_assgn76317;
    reg [31:0] z7631_assgn76318;
    reg [31:0] z3366_assgn3366;
    reg [31:0] i2_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7635_assgn7635;
    reg [31:0] z7635_assgn76350;
    reg [31:0] z7635_assgn76351;
    reg [31:0] z7635_assgn76352;
    reg [31:0] z7635_assgn76353;
    reg [31:0] z7635_assgn76354;
    reg [31:0] z7635_assgn76355;
    reg [31:0] z7635_assgn76356;
    reg [31:0] z7635_assgn76357;
    reg [31:0] z7635_assgn76358;
    reg [31:0] z3368_assgn3368;
    reg [31:0] i3_comar2_G4_mul2_G16_mul2_G256_inv0_reg;
    wire [31:0] i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0;
    reg [31:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] y1_4_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] z7657_assgn7657;
    reg [31:0] z7657_assgn76570;
    reg [31:0] z7657_assgn76571;
    reg [31:0] z7657_assgn76572;
    reg [31:0] z7657_assgn76573;
    reg [31:0] z7657_assgn76574;
    reg [31:0] z7657_assgn76575;
    reg [31:0] z7657_assgn76576;
    reg [31:0] z7657_assgn76577;
    reg [31:0] z7657_assgn76578;
    reg [31:0] z7657_assgn76579;
    reg [31:0] z7657_assgn765710;
    reg [31:0] z3387_assgn3387;
    wire [31:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [31:0] q0_0_G16_mul2_G256_inv0;
    wire [31:0] q1_0_G16_mul2_G256_inv0;
    wire [31:0] q0_G16_mul2_G256_inv0;
    wire [31:0] q1_G16_mul2_G256_inv0;
    wire [31:0] p0ls2_G16_mul2_G256_inv0;
    wire [31:0] z7671_assgn7671;
    reg [31:0] z7671_assgn76710;
    reg [31:0] z7671_assgn76711;
    reg [31:0] z7671_assgn76712;
    reg [31:0] z7671_assgn76713;
    reg [31:0] z7671_assgn76714;
    reg [31:0] z7671_assgn76715;
    reg [31:0] z7671_assgn76716;
    reg [31:0] z7671_assgn76717;
    reg [31:0] z7671_assgn76718;
    reg [31:0] z7671_assgn76719;
    reg [31:0] z7671_assgn767110;
    reg [31:0] z3399_assgn3399;
    wire [31:0] p1ls2_G16_mul2_G256_inv0;
    wire [31:0] q0_G256_inv0;
    wire [31:0] q1_G256_inv0;
    wire [31:0] p0ls4_G256_inv0;
    wire [31:0] z7681_assgn7681;
    reg [31:0] z7681_assgn76810;
    reg [31:0] z7681_assgn76811;
    reg [31:0] z7681_assgn76812;
    reg [31:0] z7681_assgn76813;
    reg [31:0] z7681_assgn76814;
    reg [31:0] z7681_assgn76815;
    reg [31:0] z7681_assgn76816;
    reg [31:0] z7681_assgn76817;
    reg [31:0] z7681_assgn76818;
    reg [31:0] z7681_assgn76819;
    reg [31:0] z7681_assgn768110;
    reg [31:0] z3407_assgn3407;
    wire [31:0] p1ls4_G256_inv0;
    wire [31:0] t4;
    wire [31:0] t5;
    wire [31:0] y_G256_newbasis1;
    wire [31:0] tempy1_G256_newbasis1;
    wire [31:0] cond1_G256_newbasis1;
    wire [31:0] negCond1_G256_newbasis1;
    wire [31:0] yxorb1_G256_newbasis1;
    wire [31:0] ny1_G256_newbasis1;
    wire [31:0] tempyIntoNegCond1_G256_newbasis1;
    wire [31:0] y1_G256_newbasis1;
    wire [31:0] x1_G256_newbasis1;
    wire [31:0] tempy2_G256_newbasis1;
    wire [31:0] cond2_G256_newbasis1;
    wire [31:0] negCond2_G256_newbasis1;
    wire [31:0] yxorb2_G256_newbasis1;
    wire [31:0] ny2_G256_newbasis1;
    wire [31:0] tempyIntoNegCond2_G256_newbasis1;
    wire [31:0] y2_G256_newbasis1;
    wire [31:0] x2_G256_newbasis1;
    wire [31:0] tempy3_G256_newbasis1;
    wire [31:0] cond3_G256_newbasis1;
    wire [31:0] negCond3_G256_newbasis1;
    wire [31:0] yxorb3_G256_newbasis1;
    wire [31:0] ny3_G256_newbasis1;
    wire [31:0] tempyIntoNegCond3_G256_newbasis1;
    wire [31:0] y3_G256_newbasis1;
    wire [31:0] x3_G256_newbasis1;
    wire [31:0] tempy4_G256_newbasis1;
    wire [31:0] cond4_G256_newbasis1;
    wire [31:0] negCond4_G256_newbasis1;
    wire [31:0] yxorb4_G256_newbasis1;
    wire [31:0] ny4_G256_newbasis1;
    wire [31:0] tempyIntoNegCond4_G256_newbasis1;
    wire [31:0] y4_G256_newbasis1;
    wire [31:0] x4_G256_newbasis1;
    wire [31:0] tempy5_G256_newbasis1;
    wire [31:0] cond5_G256_newbasis1;
    wire [31:0] negCond5_G256_newbasis1;
    wire [31:0] yxorb5_G256_newbasis1;
    wire [31:0] ny5_G256_newbasis1;
    wire [31:0] tempyIntoNegCond5_G256_newbasis1;
    wire [31:0] y5_G256_newbasis1;
    wire [31:0] x5_G256_newbasis1;
    wire [31:0] tempy6_G256_newbasis1;
    wire [31:0] cond6_G256_newbasis1;
    wire [31:0] negCond6_G256_newbasis1;
    wire [31:0] yxorb6_G256_newbasis1;
    wire [31:0] ny6_G256_newbasis1;
    wire [31:0] tempyIntoNegCond6_G256_newbasis1;
    wire [31:0] y6_G256_newbasis1;
    wire [31:0] x6_G256_newbasis1;
    wire [31:0] tempy7_G256_newbasis1;
    wire [31:0] cond7_G256_newbasis1;
    wire [31:0] negCond7_G256_newbasis1;
    wire [31:0] yxorb7_G256_newbasis1;
    wire [31:0] ny7_G256_newbasis1;
    wire [31:0] tempyIntoNegCond7_G256_newbasis1;
    wire [31:0] y7_G256_newbasis1;
    wire [31:0] x7_G256_newbasis1;
    wire [31:0] tempy8_G256_newbasis1;
    wire [31:0] cond8_G256_newbasis1;
    wire [31:0] negCond8_G256_newbasis1;
    wire [31:0] yxorb8_G256_newbasis1;
    wire [31:0] ny8_G256_newbasis1;
    wire [31:0] tempyIntoNegCond8_G256_newbasis1;
    wire [31:0] y8_G256_newbasis1;
    wire [31:0] z7817_assgn7817;
    reg [31:0] z7817_assgn78170;
    reg [31:0] z7817_assgn78171;
    reg [31:0] z7817_assgn78172;
    reg [31:0] z7817_assgn78173;
    reg [31:0] z7817_assgn78174;
    reg [31:0] z7817_assgn78175;
    reg [31:0] z7817_assgn78176;
    reg [31:0] z7817_assgn78177;
    reg [31:0] z7817_assgn78178;
    reg [31:0] z7817_assgn78179;
    reg [31:0] z7817_assgn781710;
    reg [31:0] x8_G256_newbasis1;
    wire [31:0] t6;
    wire [31:0] z_y_G256_newbasis1;
    wire [31:0] z_tempy1_G256_newbasis1;
    wire [31:0] z7825_assgn7825;
    reg [31:0] z7825_assgn78250;
    reg [31:0] z7825_assgn78251;
    reg [31:0] z7825_assgn78252;
    reg [31:0] z7825_assgn78253;
    reg [31:0] z7825_assgn78254;
    reg [31:0] z7825_assgn78255;
    reg [31:0] z7825_assgn78256;
    reg [31:0] z7825_assgn78257;
    reg [31:0] z7825_assgn78258;
    reg [31:0] z7825_assgn78259;
    reg [31:0] z7825_assgn782510;
    reg [31:0] z3549_assgn3549;
    wire [31:0] z_cond1_G256_newbasis1;
    wire [31:0] z_negCond1_G256_newbasis1;
    wire [31:0] z_yxorb1_G256_newbasis1;
    wire [31:0] z7833_assgn7833;
    reg [31:0] z7833_assgn78330;
    reg [31:0] z7833_assgn78331;
    reg [31:0] z7833_assgn78332;
    reg [31:0] z7833_assgn78333;
    reg [31:0] z7833_assgn78334;
    reg [31:0] z7833_assgn78335;
    reg [31:0] z7833_assgn78336;
    reg [31:0] z7833_assgn78337;
    reg [31:0] z7833_assgn78338;
    reg [31:0] z7833_assgn78339;
    reg [31:0] z7833_assgn783310;
    reg [31:0] z3555_assgn3555;
    wire [31:0] z_ny1_G256_newbasis1;
    wire [31:0] z7837_assgn7837;
    reg [31:0] z7837_assgn78370;
    reg [31:0] z7837_assgn78371;
    reg [31:0] z7837_assgn78372;
    reg [31:0] z7837_assgn78373;
    reg [31:0] z7837_assgn78374;
    reg [31:0] z7837_assgn78375;
    reg [31:0] z7837_assgn78376;
    reg [31:0] z7837_assgn78377;
    reg [31:0] z7837_assgn78378;
    reg [31:0] z7837_assgn78379;
    reg [31:0] z7837_assgn783710;
    reg [31:0] z3558_assgn3558;
    wire [31:0] z_tempyIntoNegCond1_G256_newbasis1;
    wire [31:0] z_y1_G256_newbasis1;
    wire [31:0] z7843_assgn7843;
    reg [31:0] z7843_assgn78430;
    reg [31:0] z7843_assgn78431;
    reg [31:0] z7843_assgn78432;
    reg [31:0] z7843_assgn78433;
    reg [31:0] z7843_assgn78434;
    reg [31:0] z7843_assgn78435;
    reg [31:0] z7843_assgn78436;
    reg [31:0] z7843_assgn78437;
    reg [31:0] z7843_assgn78438;
    reg [31:0] z7843_assgn78439;
    reg [31:0] z7843_assgn784310;
    reg [31:0] z3561_assgn3561;
    wire [31:0] z_x1_G256_newbasis1;
    wire [31:0] z_tempy2_G256_newbasis1;
    wire [31:0] z7849_assgn7849;
    reg [31:0] z7849_assgn78490;
    reg [31:0] z7849_assgn78491;
    reg [31:0] z7849_assgn78492;
    reg [31:0] z7849_assgn78493;
    reg [31:0] z7849_assgn78494;
    reg [31:0] z7849_assgn78495;
    reg [31:0] z7849_assgn78496;
    reg [31:0] z7849_assgn78497;
    reg [31:0] z7849_assgn78498;
    reg [31:0] z7849_assgn78499;
    reg [31:0] z7849_assgn784910;
    reg [31:0] z3565_assgn3565;
    wire [31:0] z_cond2_G256_newbasis1;
    wire [31:0] z_negCond2_G256_newbasis1;
    wire [31:0] z7855_assgn7855;
    reg [31:0] z7855_assgn78550;
    reg [31:0] z7855_assgn78551;
    reg [31:0] z7855_assgn78552;
    reg [31:0] z7855_assgn78553;
    reg [31:0] z7855_assgn78554;
    reg [31:0] z7855_assgn78555;
    reg [31:0] z7855_assgn78556;
    reg [31:0] z7855_assgn78557;
    reg [31:0] z7855_assgn78558;
    reg [31:0] z7855_assgn78559;
    reg [31:0] z7855_assgn785510;
    reg [31:0] z3569_assgn3569;
    wire [31:0] z_yxorb2_G256_newbasis1;
    wire [31:0] z_ny2_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond2_G256_newbasis1;
    wire [31:0] z_y2_G256_newbasis1;
    wire [31:0] z7865_assgn7865;
    reg [31:0] z7865_assgn78650;
    reg [31:0] z7865_assgn78651;
    reg [31:0] z7865_assgn78652;
    reg [31:0] z7865_assgn78653;
    reg [31:0] z7865_assgn78654;
    reg [31:0] z7865_assgn78655;
    reg [31:0] z7865_assgn78656;
    reg [31:0] z7865_assgn78657;
    reg [31:0] z7865_assgn78658;
    reg [31:0] z7865_assgn78659;
    reg [31:0] z7865_assgn786510;
    reg [31:0] z3577_assgn3577;
    wire [31:0] z_x2_G256_newbasis1;
    wire [31:0] z_tempy3_G256_newbasis1;
    wire [31:0] z7871_assgn7871;
    reg [31:0] z7871_assgn78710;
    reg [31:0] z7871_assgn78711;
    reg [31:0] z7871_assgn78712;
    reg [31:0] z7871_assgn78713;
    reg [31:0] z7871_assgn78714;
    reg [31:0] z7871_assgn78715;
    reg [31:0] z7871_assgn78716;
    reg [31:0] z7871_assgn78717;
    reg [31:0] z7871_assgn78718;
    reg [31:0] z7871_assgn78719;
    reg [31:0] z7871_assgn787110;
    reg [31:0] z3581_assgn3581;
    wire [31:0] z_cond3_G256_newbasis1;
    wire [31:0] z_negCond3_G256_newbasis1;
    wire [31:0] z7877_assgn7877;
    reg [31:0] z7877_assgn78770;
    reg [31:0] z7877_assgn78771;
    reg [31:0] z7877_assgn78772;
    reg [31:0] z7877_assgn78773;
    reg [31:0] z7877_assgn78774;
    reg [31:0] z7877_assgn78775;
    reg [31:0] z7877_assgn78776;
    reg [31:0] z7877_assgn78777;
    reg [31:0] z7877_assgn78778;
    reg [31:0] z7877_assgn78779;
    reg [31:0] z7877_assgn787710;
    reg [31:0] z3585_assgn3585;
    wire [31:0] z_yxorb3_G256_newbasis1;
    wire [31:0] z_ny3_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond3_G256_newbasis1;
    wire [31:0] z_y3_G256_newbasis1;
    wire [31:0] z7887_assgn7887;
    reg [31:0] z7887_assgn78870;
    reg [31:0] z7887_assgn78871;
    reg [31:0] z7887_assgn78872;
    reg [31:0] z7887_assgn78873;
    reg [31:0] z7887_assgn78874;
    reg [31:0] z7887_assgn78875;
    reg [31:0] z7887_assgn78876;
    reg [31:0] z7887_assgn78877;
    reg [31:0] z7887_assgn78878;
    reg [31:0] z7887_assgn78879;
    reg [31:0] z7887_assgn788710;
    reg [31:0] z3593_assgn3593;
    wire [31:0] z_x3_G256_newbasis1;
    wire [31:0] z_tempy4_G256_newbasis1;
    wire [31:0] z7893_assgn7893;
    reg [31:0] z7893_assgn78930;
    reg [31:0] z7893_assgn78931;
    reg [31:0] z7893_assgn78932;
    reg [31:0] z7893_assgn78933;
    reg [31:0] z7893_assgn78934;
    reg [31:0] z7893_assgn78935;
    reg [31:0] z7893_assgn78936;
    reg [31:0] z7893_assgn78937;
    reg [31:0] z7893_assgn78938;
    reg [31:0] z7893_assgn78939;
    reg [31:0] z7893_assgn789310;
    reg [31:0] z3597_assgn3597;
    wire [31:0] z_cond4_G256_newbasis1;
    wire [31:0] z_negCond4_G256_newbasis1;
    wire [31:0] z7899_assgn7899;
    reg [31:0] z7899_assgn78990;
    reg [31:0] z7899_assgn78991;
    reg [31:0] z7899_assgn78992;
    reg [31:0] z7899_assgn78993;
    reg [31:0] z7899_assgn78994;
    reg [31:0] z7899_assgn78995;
    reg [31:0] z7899_assgn78996;
    reg [31:0] z7899_assgn78997;
    reg [31:0] z7899_assgn78998;
    reg [31:0] z7899_assgn78999;
    reg [31:0] z7899_assgn789910;
    reg [31:0] z3601_assgn3601;
    wire [31:0] z_yxorb4_G256_newbasis1;
    wire [31:0] z_ny4_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond4_G256_newbasis1;
    wire [31:0] z_y4_G256_newbasis1;
    wire [31:0] z7909_assgn7909;
    reg [31:0] z7909_assgn79090;
    reg [31:0] z7909_assgn79091;
    reg [31:0] z7909_assgn79092;
    reg [31:0] z7909_assgn79093;
    reg [31:0] z7909_assgn79094;
    reg [31:0] z7909_assgn79095;
    reg [31:0] z7909_assgn79096;
    reg [31:0] z7909_assgn79097;
    reg [31:0] z7909_assgn79098;
    reg [31:0] z7909_assgn79099;
    reg [31:0] z7909_assgn790910;
    reg [31:0] z3609_assgn3609;
    wire [31:0] z_x4_G256_newbasis1;
    wire [31:0] z_tempy5_G256_newbasis1;
    wire [31:0] z7915_assgn7915;
    reg [31:0] z7915_assgn79150;
    reg [31:0] z7915_assgn79151;
    reg [31:0] z7915_assgn79152;
    reg [31:0] z7915_assgn79153;
    reg [31:0] z7915_assgn79154;
    reg [31:0] z7915_assgn79155;
    reg [31:0] z7915_assgn79156;
    reg [31:0] z7915_assgn79157;
    reg [31:0] z7915_assgn79158;
    reg [31:0] z7915_assgn79159;
    reg [31:0] z7915_assgn791510;
    reg [31:0] z3613_assgn3613;
    wire [31:0] z_cond5_G256_newbasis1;
    wire [31:0] z_negCond5_G256_newbasis1;
    wire [31:0] z7921_assgn7921;
    reg [31:0] z7921_assgn79210;
    reg [31:0] z7921_assgn79211;
    reg [31:0] z7921_assgn79212;
    reg [31:0] z7921_assgn79213;
    reg [31:0] z7921_assgn79214;
    reg [31:0] z7921_assgn79215;
    reg [31:0] z7921_assgn79216;
    reg [31:0] z7921_assgn79217;
    reg [31:0] z7921_assgn79218;
    reg [31:0] z7921_assgn79219;
    reg [31:0] z7921_assgn792110;
    reg [31:0] z3617_assgn3617;
    wire [31:0] z_yxorb5_G256_newbasis1;
    wire [31:0] z_ny5_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond5_G256_newbasis1;
    wire [31:0] z_y5_G256_newbasis1;
    wire [31:0] z7931_assgn7931;
    reg [31:0] z7931_assgn79310;
    reg [31:0] z7931_assgn79311;
    reg [31:0] z7931_assgn79312;
    reg [31:0] z7931_assgn79313;
    reg [31:0] z7931_assgn79314;
    reg [31:0] z7931_assgn79315;
    reg [31:0] z7931_assgn79316;
    reg [31:0] z7931_assgn79317;
    reg [31:0] z7931_assgn79318;
    reg [31:0] z7931_assgn79319;
    reg [31:0] z7931_assgn793110;
    reg [31:0] z3625_assgn3625;
    wire [31:0] z_x5_G256_newbasis1;
    wire [31:0] z_tempy6_G256_newbasis1;
    wire [31:0] z7937_assgn7937;
    reg [31:0] z7937_assgn79370;
    reg [31:0] z7937_assgn79371;
    reg [31:0] z7937_assgn79372;
    reg [31:0] z7937_assgn79373;
    reg [31:0] z7937_assgn79374;
    reg [31:0] z7937_assgn79375;
    reg [31:0] z7937_assgn79376;
    reg [31:0] z7937_assgn79377;
    reg [31:0] z7937_assgn79378;
    reg [31:0] z7937_assgn79379;
    reg [31:0] z7937_assgn793710;
    reg [31:0] z3629_assgn3629;
    wire [31:0] z_cond6_G256_newbasis1;
    wire [31:0] z_negCond6_G256_newbasis1;
    wire [31:0] z7943_assgn7943;
    reg [31:0] z7943_assgn79430;
    reg [31:0] z7943_assgn79431;
    reg [31:0] z7943_assgn79432;
    reg [31:0] z7943_assgn79433;
    reg [31:0] z7943_assgn79434;
    reg [31:0] z7943_assgn79435;
    reg [31:0] z7943_assgn79436;
    reg [31:0] z7943_assgn79437;
    reg [31:0] z7943_assgn79438;
    reg [31:0] z7943_assgn79439;
    reg [31:0] z7943_assgn794310;
    reg [31:0] z3633_assgn3633;
    wire [31:0] z_yxorb6_G256_newbasis1;
    wire [31:0] z_ny6_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond6_G256_newbasis1;
    wire [31:0] z_y6_G256_newbasis1;
    wire [31:0] z7953_assgn7953;
    reg [31:0] z7953_assgn79530;
    reg [31:0] z7953_assgn79531;
    reg [31:0] z7953_assgn79532;
    reg [31:0] z7953_assgn79533;
    reg [31:0] z7953_assgn79534;
    reg [31:0] z7953_assgn79535;
    reg [31:0] z7953_assgn79536;
    reg [31:0] z7953_assgn79537;
    reg [31:0] z7953_assgn79538;
    reg [31:0] z7953_assgn79539;
    reg [31:0] z7953_assgn795310;
    reg [31:0] z3641_assgn3641;
    wire [31:0] z_x6_G256_newbasis1;
    wire [31:0] z_tempy7_G256_newbasis1;
    wire [31:0] z7959_assgn7959;
    reg [31:0] z7959_assgn79590;
    reg [31:0] z7959_assgn79591;
    reg [31:0] z7959_assgn79592;
    reg [31:0] z7959_assgn79593;
    reg [31:0] z7959_assgn79594;
    reg [31:0] z7959_assgn79595;
    reg [31:0] z7959_assgn79596;
    reg [31:0] z7959_assgn79597;
    reg [31:0] z7959_assgn79598;
    reg [31:0] z7959_assgn79599;
    reg [31:0] z7959_assgn795910;
    reg [31:0] z3645_assgn3645;
    wire [31:0] z_cond7_G256_newbasis1;
    wire [31:0] z_negCond7_G256_newbasis1;
    wire [31:0] z7965_assgn7965;
    reg [31:0] z7965_assgn79650;
    reg [31:0] z7965_assgn79651;
    reg [31:0] z7965_assgn79652;
    reg [31:0] z7965_assgn79653;
    reg [31:0] z7965_assgn79654;
    reg [31:0] z7965_assgn79655;
    reg [31:0] z7965_assgn79656;
    reg [31:0] z7965_assgn79657;
    reg [31:0] z7965_assgn79658;
    reg [31:0] z7965_assgn79659;
    reg [31:0] z7965_assgn796510;
    reg [31:0] z3649_assgn3649;
    wire [31:0] z_yxorb7_G256_newbasis1;
    wire [31:0] z_ny7_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond7_G256_newbasis1;
    wire [31:0] z_y7_G256_newbasis1;
    wire [31:0] z7975_assgn7975;
    reg [31:0] z7975_assgn79750;
    reg [31:0] z7975_assgn79751;
    reg [31:0] z7975_assgn79752;
    reg [31:0] z7975_assgn79753;
    reg [31:0] z7975_assgn79754;
    reg [31:0] z7975_assgn79755;
    reg [31:0] z7975_assgn79756;
    reg [31:0] z7975_assgn79757;
    reg [31:0] z7975_assgn79758;
    reg [31:0] z7975_assgn79759;
    reg [31:0] z7975_assgn797510;
    reg [31:0] z3657_assgn3657;
    wire [31:0] z_x7_G256_newbasis1;
    wire [31:0] z_tempy8_G256_newbasis1;
    wire [31:0] z7981_assgn7981;
    reg [31:0] z7981_assgn79810;
    reg [31:0] z7981_assgn79811;
    reg [31:0] z7981_assgn79812;
    reg [31:0] z7981_assgn79813;
    reg [31:0] z7981_assgn79814;
    reg [31:0] z7981_assgn79815;
    reg [31:0] z7981_assgn79816;
    reg [31:0] z7981_assgn79817;
    reg [31:0] z7981_assgn79818;
    reg [31:0] z7981_assgn79819;
    reg [31:0] z7981_assgn798110;
    reg [31:0] z3661_assgn3661;
    wire [31:0] z_cond8_G256_newbasis1;
    wire [31:0] z_negCond8_G256_newbasis1;
    wire [31:0] z7987_assgn7987;
    reg [31:0] z7987_assgn79870;
    reg [31:0] z7987_assgn79871;
    reg [31:0] z7987_assgn79872;
    reg [31:0] z7987_assgn79873;
    reg [31:0] z7987_assgn79874;
    reg [31:0] z7987_assgn79875;
    reg [31:0] z7987_assgn79876;
    reg [31:0] z7987_assgn79877;
    reg [31:0] z7987_assgn79878;
    reg [31:0] z7987_assgn79879;
    reg [31:0] z7987_assgn798710;
    reg [31:0] z3665_assgn3665;
    wire [31:0] z_yxorb8_G256_newbasis1;
    wire [31:0] z_ny8_G256_newbasis1;
    wire [31:0] z_tempyIntoNegCond8_G256_newbasis1;
    wire [31:0] z_y8_G256_newbasis1;
    wire [31:0] z7997_assgn7997;
    reg [31:0] z7997_assgn79970;
    reg [31:0] z7997_assgn79971;
    reg [31:0] z7997_assgn79972;
    reg [31:0] z7997_assgn79973;
    reg [31:0] z7997_assgn79974;
    reg [31:0] z7997_assgn79975;
    reg [31:0] z7997_assgn79976;
    reg [31:0] z7997_assgn79977;
    reg [31:0] z7997_assgn79978;
    reg [31:0] z7997_assgn79979;
    reg [31:0] z7997_assgn799710;
    reg [31:0] z3673_assgn3673;
    wire [31:0] z_x8_G256_newbasis1;
    wire [31:0] t7;
    wire [31:0] z8003_assgn8003;
    reg [31:0] z8003_assgn80030;
    reg [31:0] z8003_assgn80031;
    reg [31:0] z8003_assgn80032;
    reg [31:0] z8003_assgn80033;
    reg [31:0] z8003_assgn80034;
    reg [31:0] z8003_assgn80035;
    reg [31:0] z8003_assgn80036;
    reg [31:0] z8003_assgn80037;
    reg [31:0] z8003_assgn80038;
    reg [31:0] z8003_assgn80039;
    reg [31:0] z8003_assgn800310;

    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempyIntoNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempyIntoNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempyIntoNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempyIntoNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempyIntoNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempyIntoNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempyIntoNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempyIntoNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempyIntoNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempyIntoNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempyIntoNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempyIntoNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempyIntoNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempyIntoNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempyIntoNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempyIntoNegCond8_G256_newbasis0);
    assign z3873_assgn3873 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempyIntoNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempyIntoNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempyIntoNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempyIntoNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempyIntoNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempyIntoNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempyIntoNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempyIntoNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempyIntoNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempyIntoNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempyIntoNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempyIntoNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempyIntoNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempyIntoNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempyIntoNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempyIntoNegCond8_G256_newbasis0);
    assign z4005_assgn4005 = (z_x7_G256_newbasis0 >> dec_1_inp);
    assign t3 = z_y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a1_0_G256_inv0 = (t3 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a1xorb1_G256_inv0 = (a1_G256_inv0 ^ b1_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul0_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ d1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul0_G16_mul0_G256_inv0 = (m0_comar0_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_comar0_G4_mul0_G16_mul0_G256_inv0 = (m3_comar0_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_comar0_G4_mul0_G16_mul0_G256_inv0 = (m0_comar0_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_comar0_G4_mul0_G16_mul0_G256_inv0 = (m3_comar0_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0_comar0_G4_mul0_G16_mul0_G256_inv0 = (p1_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_comar0_G4_mul0_G16_mul0_G256_inv0 = (p2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_comar0_G4_mul0_G16_mul0_G256_inv0 = (p3_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i3_comar0_G4_mul0_G16_mul0_G256_inv0 = (p4_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0 = (i1_comar0_G4_mul0_G16_mul0_G256_inv0_reg ^ i2_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0 = (i0_comar0_G4_mul0_G16_mul0_G256_inv0_reg ^ i3_comar0_G4_mul0_G16_mul0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul0_G16_mul0_G256_inv0 = (r00_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul0_G16_mul0_G256_inv0 = (m0_comar1_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_comar1_G4_mul0_G16_mul0_G256_inv0 = (m3_comar1_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_comar1_G4_mul0_G16_mul0_G256_inv0 = (m0_comar1_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_comar1_G4_mul0_G16_mul0_G256_inv0 = (m3_comar1_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0_comar1_G4_mul0_G16_mul0_G256_inv0 = (p1_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_comar1_G4_mul0_G16_mul0_G256_inv0 = (p2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_comar1_G4_mul0_G16_mul0_G256_inv0 = (p3_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i3_comar1_G4_mul0_G16_mul0_G256_inv0 = (p4_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0 = (i1_comar1_G4_mul0_G16_mul0_G256_inv0_reg ^ i2_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0 = (i0_comar1_G4_mul0_G16_mul0_G256_inv0_reg ^ i3_comar1_G4_mul0_G16_mul0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul0_G16_mul0_G256_inv0 = (r00_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul0_G256_inv0 = (d1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul0_G256_inv0 = (d0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul0_G16_mul0_G256_inv0 = (m0_comar2_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p3_comar2_G4_mul0_G16_mul0_G256_inv0 = (m3_comar2_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p1_comar2_G4_mul0_G16_mul0_G256_inv0 = (m0_comar2_G4_mul0_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign p4_comar2_G4_mul0_G16_mul0_G256_inv0 = (m3_comar2_G4_mul0_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0_comar2_G4_mul0_G16_mul0_G256_inv0 = (p1_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1_comar2_G4_mul0_G16_mul0_G256_inv0 = (p2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i2_comar2_G4_mul0_G16_mul0_G256_inv0 = (p3_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i3_comar2_G4_mul0_G16_mul0_G256_inv0 = (p4_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0 = (i1_comar2_G4_mul0_G16_mul0_G256_inv0_reg ^ i2_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0 = (i0_comar2_G4_mul0_G16_mul0_G256_inv0_reg ^ i3_comar2_G4_mul0_G16_mul0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul0_G16_mul0_G256_inv0 = (r00_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp);
    assign z4371_assgn4371 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << z691_assgn691);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_2_inp);
    assign z4381_assgn4381 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z699_assgn699);
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign z4387_assgn4387 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> z703_assgn703);
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_1_inp);
    assign z4393_assgn4393 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & z707_assgn707);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign z4405_assgn4405 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << z717_assgn717);
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ d1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul0_G256_inv0 = (cxord_1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul0_G256_inv0 = (cxord_0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul1_G16_mul0_G256_inv0 = (m0_comar0_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_comar0_G4_mul1_G16_mul0_G256_inv0 = (m3_comar0_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_comar0_G4_mul1_G16_mul0_G256_inv0 = (m0_comar0_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_comar0_G4_mul1_G16_mul0_G256_inv0 = (m3_comar0_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0_comar0_G4_mul1_G16_mul0_G256_inv0 = (p1_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_comar0_G4_mul1_G16_mul0_G256_inv0 = (p2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_comar0_G4_mul1_G16_mul0_G256_inv0 = (p3_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i3_comar0_G4_mul1_G16_mul0_G256_inv0 = (p4_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0 = (i1_comar0_G4_mul1_G16_mul0_G256_inv0_reg ^ i2_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0 = (i0_comar0_G4_mul1_G16_mul0_G256_inv0_reg ^ i3_comar0_G4_mul1_G16_mul0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul1_G16_mul0_G256_inv0 = (r00_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul1_G16_mul0_G256_inv0 = (m0_comar1_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_comar1_G4_mul1_G16_mul0_G256_inv0 = (m3_comar1_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_comar1_G4_mul1_G16_mul0_G256_inv0 = (m0_comar1_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_comar1_G4_mul1_G16_mul0_G256_inv0 = (m3_comar1_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0_comar1_G4_mul1_G16_mul0_G256_inv0 = (p1_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_comar1_G4_mul1_G16_mul0_G256_inv0 = (p2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_comar1_G4_mul1_G16_mul0_G256_inv0 = (p3_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i3_comar1_G4_mul1_G16_mul0_G256_inv0 = (p4_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0 = (i1_comar1_G4_mul1_G16_mul0_G256_inv0_reg ^ i2_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0 = (i0_comar1_G4_mul1_G16_mul0_G256_inv0_reg ^ i3_comar1_G4_mul1_G16_mul0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul1_G16_mul0_G256_inv0 = (r00_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul0_G256_inv0 = (d1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul0_G256_inv0 = (d0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul1_G16_mul0_G256_inv0 = (m0_comar2_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p3_comar2_G4_mul1_G16_mul0_G256_inv0 = (m3_comar2_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p1_comar2_G4_mul1_G16_mul0_G256_inv0 = (m0_comar2_G4_mul1_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign p4_comar2_G4_mul1_G16_mul0_G256_inv0 = (m3_comar2_G4_mul1_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0_comar2_G4_mul1_G16_mul0_G256_inv0 = (p1_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1_comar2_G4_mul1_G16_mul0_G256_inv0 = (p2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i2_comar2_G4_mul1_G16_mul0_G256_inv0 = (p3_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i3_comar2_G4_mul1_G16_mul0_G256_inv0 = (p4_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0 = (i1_comar2_G4_mul1_G16_mul0_G256_inv0_reg ^ i2_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0 = (i0_comar2_G4_mul1_G16_mul0_G256_inv0_reg ^ i3_comar2_G4_mul1_G16_mul0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul1_G16_mul0_G256_inv0 = (r00_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp);
    assign z4625_assgn4625 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << z935_assgn935);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ d1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul0_G256_inv0 = (cxord_1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul0_G256_inv0 = (cxord_0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul2_G16_mul0_G256_inv0 = (m0_comar0_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_comar0_G4_mul2_G16_mul0_G256_inv0 = (m3_comar0_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_comar0_G4_mul2_G16_mul0_G256_inv0 = (m0_comar0_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_comar0_G4_mul2_G16_mul0_G256_inv0 = (m3_comar0_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0_comar0_G4_mul2_G16_mul0_G256_inv0 = (p1_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_comar0_G4_mul2_G16_mul0_G256_inv0 = (p2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_comar0_G4_mul2_G16_mul0_G256_inv0 = (p3_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i3_comar0_G4_mul2_G16_mul0_G256_inv0 = (p4_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0 = (i1_comar0_G4_mul2_G16_mul0_G256_inv0_reg ^ i2_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0 = (i0_comar0_G4_mul2_G16_mul0_G256_inv0_reg ^ i3_comar0_G4_mul2_G16_mul0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul2_G16_mul0_G256_inv0 = (r00_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul2_G16_mul0_G256_inv0 = (m0_comar1_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_comar1_G4_mul2_G16_mul0_G256_inv0 = (m3_comar1_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_comar1_G4_mul2_G16_mul0_G256_inv0 = (m0_comar1_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_comar1_G4_mul2_G16_mul0_G256_inv0 = (m3_comar1_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0_comar1_G4_mul2_G16_mul0_G256_inv0 = (p1_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_comar1_G4_mul2_G16_mul0_G256_inv0 = (p2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_comar1_G4_mul2_G16_mul0_G256_inv0 = (p3_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i3_comar1_G4_mul2_G16_mul0_G256_inv0 = (p4_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0 = (i1_comar1_G4_mul2_G16_mul0_G256_inv0_reg ^ i2_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0 = (i0_comar1_G4_mul2_G16_mul0_G256_inv0_reg ^ i3_comar1_G4_mul2_G16_mul0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul2_G16_mul0_G256_inv0 = (r00_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul0_G256_inv0 = (d1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul0_G256_inv0 = (d0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul2_G16_mul0_G256_inv0 = (m0_comar2_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p3_comar2_G4_mul2_G16_mul0_G256_inv0 = (m3_comar2_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p1_comar2_G4_mul2_G16_mul0_G256_inv0 = (m0_comar2_G4_mul2_G16_mul0_G256_inv0_reg & m2_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign p4_comar2_G4_mul2_G16_mul0_G256_inv0 = (m3_comar2_G4_mul2_G16_mul0_G256_inv0_reg & m1_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0_comar2_G4_mul2_G16_mul0_G256_inv0 = (p1_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1_comar2_G4_mul2_G16_mul0_G256_inv0 = (p2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i2_comar2_G4_mul2_G16_mul0_G256_inv0 = (p3_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i3_comar2_G4_mul2_G16_mul0_G256_inv0 = (p4_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0 = (i1_comar2_G4_mul2_G16_mul0_G256_inv0_reg ^ i2_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0 = (i0_comar2_G4_mul2_G16_mul0_G256_inv0_reg ^ i3_comar2_G4_mul2_G16_mul0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul2_G16_mul0_G256_inv0 = (r00_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp);
    assign z4847_assgn4847 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << z1155_assgn1155);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << dec_2_inp);
    assign z4861_assgn4861 = dec_2_inp;
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << z1167_assgn1167);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign c0xord0_G256_inv0 = (c0_G256_inv0 ^ d0_G256_inv0);
    assign z4871_assgn4871 = c1_G256_inv0;
    assign c1xord1_G256_inv0 = (z1176_assgn1176 ^ d1_G256_inv0);
    assign r00_G16_inv0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_inv0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_inv0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_inv0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_inv0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_inv0_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_12_inp);
    assign z4889_assgn4889 = dec_12_inp;
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1191_assgn1191);
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> dec_2_inp);
    assign z4895_assgn4895 = dec_2_inp;
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> z1195_assgn1195);
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_3_inp);
    assign z4901_assgn4901 = dec_3_inp;
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & z1199_assgn1199);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a1xorb1_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 ^ b1_G16_inv0_G256_inv0);
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z4911_assgn4911 = dec_2_inp;
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1207_assgn1207);
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z4917_assgn4917 = dec_1_inp;
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> z1211_assgn1211);
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z4923_assgn4923 = dec_1_inp;
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & z1215_assgn1215);
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp);
    assign z4929_assgn4929 = dec_1_inp;
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << z1219_assgn1219);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z4939_assgn4939 = dec_2_inp;
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1227_assgn1227);
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z4945_assgn4945 = dec_1_inp;
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> z1231_assgn1231);
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z4951_assgn4951 = dec_1_inp;
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & z1235_assgn1235);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign z4963_assgn4963 = dec_1_inp;
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << z1245_assgn1245);
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul3_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul3_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul3_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z4987_assgn4987 = dec_2_inp;
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1267_assgn1267);
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z4993_assgn4993 = dec_1_inp;
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> z1271_assgn1271);
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z4999_assgn4999 = dec_1_inp;
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1275_assgn1275);
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5005_assgn5005 = dec_2_inp;
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1279_assgn1279);
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5011_assgn5011 = dec_1_inp;
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> z1283_assgn1283);
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5017_assgn5017 = dec_1_inp;
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1287_assgn1287);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ d1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign z5043_assgn5043 = r10_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign m1_comar0_G4_mul3_G16_inv0_G256_inv0 = (cxord_1_G4_mul3_G16_inv0_G256_inv0 ^ z1311_assgn1311);
    assign m2_comar0_G4_mul3_G16_inv0_G256_inv0 = (cxord_0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign z5049_assgn5049 = r00_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign m3_comar0_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 ^ z1315_assgn1315);
    assign z5053_assgn5053 = m0_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign p2_comar0_G4_mul3_G16_inv0_G256_inv0 = (z1318_assgn1318 & m1_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5057_assgn5057 = m2_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign p3_comar0_G4_mul3_G16_inv0_G256_inv0 = (m3_comar0_G4_mul3_G16_inv0_G256_inv0_reg & z1319_assgn1319);
    assign p1_comar0_G4_mul3_G16_inv0_G256_inv0 = (m0_comar0_G4_mul3_G16_inv0_G256_inv0_reg & m2_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_comar0_G4_mul3_G16_inv0_G256_inv0 = (m3_comar0_G4_mul3_G16_inv0_G256_inv0_reg & m1_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign i0_comar0_G4_mul3_G16_inv0_G256_inv0 = (p1_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5067_assgn5067 = r1_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign i1_comar0_G4_mul3_G16_inv0_G256_inv0 = (p2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ z1327_assgn1327);
    assign z5071_assgn5071 = r2_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign i2_comar0_G4_mul3_G16_inv0_G256_inv0 = (p3_comar0_G4_mul3_G16_inv0_G256_inv0 ^ z1329_assgn1329);
    assign z5075_assgn5075 = r3_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign i3_comar0_G4_mul3_G16_inv0_G256_inv0 = (p4_comar0_G4_mul3_G16_inv0_G256_inv0 ^ z1331_assgn1331);
    assign i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0 = (i1_comar0_G4_mul3_G16_inv0_G256_inv0_reg ^ i2_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5081_assgn5081 = i0_comar0_G4_mul3_G16_inv0_G256_inv0;
    assign i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0 = (z1336_assgn1336 ^ i3_comar0_G4_mul3_G16_inv0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul3_G16_inv0_G256_inv0 = (r00_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign z5111_assgn5111 = r10_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign m1_comar1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ z1363_assgn1363);
    assign m2_comar1_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign z5117_assgn5117 = r00_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign m3_comar1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ z1367_assgn1367);
    assign z5121_assgn5121 = m0_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign p2_comar1_G4_mul3_G16_inv0_G256_inv0 = (z1370_assgn1370 & m1_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5125_assgn5125 = m2_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign p3_comar1_G4_mul3_G16_inv0_G256_inv0 = (m3_comar1_G4_mul3_G16_inv0_G256_inv0_reg & z1371_assgn1371);
    assign p1_comar1_G4_mul3_G16_inv0_G256_inv0 = (m0_comar1_G4_mul3_G16_inv0_G256_inv0_reg & m2_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_comar1_G4_mul3_G16_inv0_G256_inv0 = (m3_comar1_G4_mul3_G16_inv0_G256_inv0_reg & m1_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign i0_comar1_G4_mul3_G16_inv0_G256_inv0 = (p1_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5135_assgn5135 = r1_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign i1_comar1_G4_mul3_G16_inv0_G256_inv0 = (p2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ z1379_assgn1379);
    assign z5139_assgn5139 = r2_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign i2_comar1_G4_mul3_G16_inv0_G256_inv0 = (p3_comar1_G4_mul3_G16_inv0_G256_inv0 ^ z1381_assgn1381);
    assign z5143_assgn5143 = r3_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign i3_comar1_G4_mul3_G16_inv0_G256_inv0 = (p4_comar1_G4_mul3_G16_inv0_G256_inv0 ^ z1383_assgn1383);
    assign i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0 = (i1_comar1_G4_mul3_G16_inv0_G256_inv0_reg ^ i2_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5149_assgn5149 = i0_comar1_G4_mul3_G16_inv0_G256_inv0;
    assign i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0 = (z1388_assgn1388 ^ i3_comar1_G4_mul3_G16_inv0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul3_G16_inv0_G256_inv0 = (r00_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign z5183_assgn5183 = r10_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign m1_comar2_G4_mul3_G16_inv0_G256_inv0 = (d1_G4_mul3_G16_inv0_G256_inv0 ^ z1419_assgn1419);
    assign m2_comar2_G4_mul3_G16_inv0_G256_inv0 = (d0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign z5189_assgn5189 = r00_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign m3_comar2_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 ^ z1423_assgn1423);
    assign z5193_assgn5193 = m0_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign p2_comar2_G4_mul3_G16_inv0_G256_inv0 = (z1426_assgn1426 & m1_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5197_assgn5197 = m2_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign p3_comar2_G4_mul3_G16_inv0_G256_inv0 = (m3_comar2_G4_mul3_G16_inv0_G256_inv0_reg & z1427_assgn1427);
    assign p1_comar2_G4_mul3_G16_inv0_G256_inv0 = (m0_comar2_G4_mul3_G16_inv0_G256_inv0_reg & m2_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign p4_comar2_G4_mul3_G16_inv0_G256_inv0 = (m3_comar2_G4_mul3_G16_inv0_G256_inv0_reg & m1_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign i0_comar2_G4_mul3_G16_inv0_G256_inv0 = (p1_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5207_assgn5207 = r1_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign i1_comar2_G4_mul3_G16_inv0_G256_inv0 = (p2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ z1435_assgn1435);
    assign z5211_assgn5211 = r2_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign i2_comar2_G4_mul3_G16_inv0_G256_inv0 = (p3_comar2_G4_mul3_G16_inv0_G256_inv0 ^ z1437_assgn1437);
    assign z5215_assgn5215 = r3_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign i3_comar2_G4_mul3_G16_inv0_G256_inv0 = (p4_comar2_G4_mul3_G16_inv0_G256_inv0 ^ z1439_assgn1439);
    assign i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0 = (i1_comar2_G4_mul3_G16_inv0_G256_inv0_reg ^ i2_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign z5221_assgn5221 = i0_comar2_G4_mul3_G16_inv0_G256_inv0;
    assign i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0 = (z1444_assgn1444 ^ i3_comar2_G4_mul3_G16_inv0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul3_G16_inv0_G256_inv0 = (r00_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << dec_1_inp);
    assign z5243_assgn5243 = dec_1_inp;
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << z1463_assgn1463);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign c0xord0_G16_inv0_G256_inv0 = (c0_G16_inv0_G256_inv0 ^ d0_G16_inv0_G256_inv0);
    assign z5253_assgn5253 = c1_G16_inv0_G256_inv0;
    assign c1xord1_G16_inv0_G256_inv0 = (z1472_assgn1472 ^ d1_G16_inv0_G256_inv0);
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5259_assgn5259 = dec_2_inp;
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1475_assgn1475);
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5265_assgn5265 = dec_1_inp;
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> z1479_assgn1479);
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5271_assgn5271 = dec_1_inp;
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & z1483_assgn1483);
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << dec_1_inp);
    assign z5277_assgn5277 = dec_1_inp;
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << z1487_assgn1487);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul4_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul4_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul4_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5299_assgn5299 = dec_2_inp;
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1507_assgn1507);
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5305_assgn5305 = dec_1_inp;
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> z1511_assgn1511);
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5311_assgn5311 = dec_1_inp;
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1515_assgn1515);
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5317_assgn5317 = dec_2_inp;
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1519_assgn1519);
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5323_assgn5323 = dec_1_inp;
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> z1523_assgn1523);
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5329_assgn5329 = dec_1_inp;
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & z1527_assgn1527);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ d1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign z5355_assgn5355 = r10_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign m1_comar0_G4_mul4_G16_inv0_G256_inv0 = (cxord_1_G4_mul4_G16_inv0_G256_inv0 ^ z1551_assgn1551);
    assign m2_comar0_G4_mul4_G16_inv0_G256_inv0 = (cxord_0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign z5361_assgn5361 = r00_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign m3_comar0_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 ^ z1555_assgn1555);
    assign z5365_assgn5365 = m0_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign p2_comar0_G4_mul4_G16_inv0_G256_inv0 = (z1558_assgn1558 & m1_comar0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5369_assgn5369 = m2_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign p3_comar0_G4_mul4_G16_inv0_G256_inv0 = (m3_comar0_G4_mul4_G16_inv0_G256_inv0_reg & z1559_assgn1559);
    assign p1_comar0_G4_mul4_G16_inv0_G256_inv0 = (m0_comar0_G4_mul4_G16_inv0_G256_inv0_reg & m2_comar0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5375_assgn5375 = m1_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign p4_comar0_G4_mul4_G16_inv0_G256_inv0 = (m3_comar0_G4_mul4_G16_inv0_G256_inv0_reg & z1563_assgn1563);
    assign i0_comar0_G4_mul4_G16_inv0_G256_inv0 = (p1_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5381_assgn5381 = r1_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign i1_comar0_G4_mul4_G16_inv0_G256_inv0 = (p2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ z1567_assgn1567);
    assign z5385_assgn5385 = r2_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign i2_comar0_G4_mul4_G16_inv0_G256_inv0 = (p3_comar0_G4_mul4_G16_inv0_G256_inv0 ^ z1569_assgn1569);
    assign z5389_assgn5389 = r3_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign i3_comar0_G4_mul4_G16_inv0_G256_inv0 = (p4_comar0_G4_mul4_G16_inv0_G256_inv0 ^ z1571_assgn1571);
    assign z5393_assgn5393 = i1_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0 = (z1574_assgn1574 ^ i2_comar0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5397_assgn5397 = i0_comar0_G4_mul4_G16_inv0_G256_inv0;
    assign i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0 = (z1576_assgn1576 ^ i3_comar0_G4_mul4_G16_inv0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul4_G16_inv0_G256_inv0 = (r00_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign z5427_assgn5427 = r10_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign m1_comar1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ z1603_assgn1603);
    assign m2_comar1_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign z5433_assgn5433 = r00_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign m3_comar1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ z1607_assgn1607);
    assign z5437_assgn5437 = m0_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign p2_comar1_G4_mul4_G16_inv0_G256_inv0 = (z1610_assgn1610 & m1_comar1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5441_assgn5441 = m2_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign p3_comar1_G4_mul4_G16_inv0_G256_inv0 = (m3_comar1_G4_mul4_G16_inv0_G256_inv0_reg & z1611_assgn1611);
    assign p1_comar1_G4_mul4_G16_inv0_G256_inv0 = (m0_comar1_G4_mul4_G16_inv0_G256_inv0_reg & m2_comar1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5447_assgn5447 = m1_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign p4_comar1_G4_mul4_G16_inv0_G256_inv0 = (m3_comar1_G4_mul4_G16_inv0_G256_inv0_reg & z1615_assgn1615);
    assign i0_comar1_G4_mul4_G16_inv0_G256_inv0 = (p1_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5453_assgn5453 = r1_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign i1_comar1_G4_mul4_G16_inv0_G256_inv0 = (p2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ z1619_assgn1619);
    assign z5457_assgn5457 = r2_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign i2_comar1_G4_mul4_G16_inv0_G256_inv0 = (p3_comar1_G4_mul4_G16_inv0_G256_inv0 ^ z1621_assgn1621);
    assign z5461_assgn5461 = r3_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign i3_comar1_G4_mul4_G16_inv0_G256_inv0 = (p4_comar1_G4_mul4_G16_inv0_G256_inv0 ^ z1623_assgn1623);
    assign z5465_assgn5465 = i1_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0 = (z1626_assgn1626 ^ i2_comar1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5469_assgn5469 = i0_comar1_G4_mul4_G16_inv0_G256_inv0;
    assign i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0 = (z1628_assgn1628 ^ i3_comar1_G4_mul4_G16_inv0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul4_G16_inv0_G256_inv0 = (r00_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign z5503_assgn5503 = r10_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign m1_comar2_G4_mul4_G16_inv0_G256_inv0 = (d1_G4_mul4_G16_inv0_G256_inv0 ^ z1659_assgn1659);
    assign m2_comar2_G4_mul4_G16_inv0_G256_inv0 = (d0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign z5509_assgn5509 = r00_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign m3_comar2_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 ^ z1663_assgn1663);
    assign z5513_assgn5513 = m0_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign p2_comar2_G4_mul4_G16_inv0_G256_inv0 = (z1666_assgn1666 & m1_comar2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5517_assgn5517 = m2_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign p3_comar2_G4_mul4_G16_inv0_G256_inv0 = (m3_comar2_G4_mul4_G16_inv0_G256_inv0_reg & z1667_assgn1667);
    assign p1_comar2_G4_mul4_G16_inv0_G256_inv0 = (m0_comar2_G4_mul4_G16_inv0_G256_inv0_reg & m2_comar2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5523_assgn5523 = m1_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign p4_comar2_G4_mul4_G16_inv0_G256_inv0 = (m3_comar2_G4_mul4_G16_inv0_G256_inv0_reg & z1671_assgn1671);
    assign i0_comar2_G4_mul4_G16_inv0_G256_inv0 = (p1_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5529_assgn5529 = r1_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign i1_comar2_G4_mul4_G16_inv0_G256_inv0 = (p2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ z1675_assgn1675);
    assign z5533_assgn5533 = r2_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign i2_comar2_G4_mul4_G16_inv0_G256_inv0 = (p3_comar2_G4_mul4_G16_inv0_G256_inv0 ^ z1677_assgn1677);
    assign z5537_assgn5537 = r3_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign i3_comar2_G4_mul4_G16_inv0_G256_inv0 = (p4_comar2_G4_mul4_G16_inv0_G256_inv0 ^ z1679_assgn1679);
    assign z5541_assgn5541 = i1_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0 = (z1682_assgn1682 ^ i2_comar2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign z5545_assgn5545 = i0_comar2_G4_mul4_G16_inv0_G256_inv0;
    assign i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0 = (z1684_assgn1684 ^ i3_comar2_G4_mul4_G16_inv0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul4_G16_inv0_G256_inv0 = (r00_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << dec_1_inp);
    assign z5567_assgn5567 = dec_1_inp;
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << z1703_assgn1703);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul5_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul5_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul5_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5589_assgn5589 = dec_2_inp;
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1723_assgn1723);
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5595_assgn5595 = dec_1_inp;
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> z1727_assgn1727);
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5601_assgn5601 = dec_1_inp;
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & z1731_assgn1731);
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign z5607_assgn5607 = dec_2_inp;
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1735_assgn1735);
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign z5613_assgn5613 = dec_1_inp;
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> z1739_assgn1739);
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign z5619_assgn5619 = dec_1_inp;
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & z1743_assgn1743);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ d1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign z5645_assgn5645 = r10_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign m1_comar0_G4_mul5_G16_inv0_G256_inv0 = (cxord_1_G4_mul5_G16_inv0_G256_inv0 ^ z1767_assgn1767);
    assign m2_comar0_G4_mul5_G16_inv0_G256_inv0 = (cxord_0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign z5651_assgn5651 = r00_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign m3_comar0_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 ^ z1771_assgn1771);
    assign z5655_assgn5655 = m0_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign p2_comar0_G4_mul5_G16_inv0_G256_inv0 = (z1774_assgn1774 & m1_comar0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5659_assgn5659 = m2_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign p3_comar0_G4_mul5_G16_inv0_G256_inv0 = (m3_comar0_G4_mul5_G16_inv0_G256_inv0_reg & z1775_assgn1775);
    assign p1_comar0_G4_mul5_G16_inv0_G256_inv0 = (m0_comar0_G4_mul5_G16_inv0_G256_inv0_reg & m2_comar0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5665_assgn5665 = m1_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign p4_comar0_G4_mul5_G16_inv0_G256_inv0 = (m3_comar0_G4_mul5_G16_inv0_G256_inv0_reg & z1779_assgn1779);
    assign i0_comar0_G4_mul5_G16_inv0_G256_inv0 = (p1_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5671_assgn5671 = r1_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign i1_comar0_G4_mul5_G16_inv0_G256_inv0 = (p2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ z1783_assgn1783);
    assign z5675_assgn5675 = r2_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign i2_comar0_G4_mul5_G16_inv0_G256_inv0 = (p3_comar0_G4_mul5_G16_inv0_G256_inv0 ^ z1785_assgn1785);
    assign z5679_assgn5679 = r3_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign i3_comar0_G4_mul5_G16_inv0_G256_inv0 = (p4_comar0_G4_mul5_G16_inv0_G256_inv0 ^ z1787_assgn1787);
    assign z5683_assgn5683 = i1_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0 = (z1790_assgn1790 ^ i2_comar0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5687_assgn5687 = i0_comar0_G4_mul5_G16_inv0_G256_inv0;
    assign i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0 = (z1792_assgn1792 ^ i3_comar0_G4_mul5_G16_inv0_G256_inv0_reg);
    assign y1_1_comar0_G4_mul5_G16_inv0_G256_inv0 = (r00_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign z5717_assgn5717 = r10_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign m1_comar1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ z1819_assgn1819);
    assign m2_comar1_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign z5723_assgn5723 = r00_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign m3_comar1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ z1823_assgn1823);
    assign z5727_assgn5727 = m0_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign p2_comar1_G4_mul5_G16_inv0_G256_inv0 = (z1826_assgn1826 & m1_comar1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5731_assgn5731 = m2_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign p3_comar1_G4_mul5_G16_inv0_G256_inv0 = (m3_comar1_G4_mul5_G16_inv0_G256_inv0_reg & z1827_assgn1827);
    assign p1_comar1_G4_mul5_G16_inv0_G256_inv0 = (m0_comar1_G4_mul5_G16_inv0_G256_inv0_reg & m2_comar1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5737_assgn5737 = m1_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign p4_comar1_G4_mul5_G16_inv0_G256_inv0 = (m3_comar1_G4_mul5_G16_inv0_G256_inv0_reg & z1831_assgn1831);
    assign i0_comar1_G4_mul5_G16_inv0_G256_inv0 = (p1_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5743_assgn5743 = r1_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign i1_comar1_G4_mul5_G16_inv0_G256_inv0 = (p2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ z1835_assgn1835);
    assign z5747_assgn5747 = r2_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign i2_comar1_G4_mul5_G16_inv0_G256_inv0 = (p3_comar1_G4_mul5_G16_inv0_G256_inv0 ^ z1837_assgn1837);
    assign z5751_assgn5751 = r3_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign i3_comar1_G4_mul5_G16_inv0_G256_inv0 = (p4_comar1_G4_mul5_G16_inv0_G256_inv0 ^ z1839_assgn1839);
    assign z5755_assgn5755 = i1_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0 = (z1842_assgn1842 ^ i2_comar1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5759_assgn5759 = i0_comar1_G4_mul5_G16_inv0_G256_inv0;
    assign i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0 = (z1844_assgn1844 ^ i3_comar1_G4_mul5_G16_inv0_G256_inv0_reg);
    assign y1_1_comar1_G4_mul5_G16_inv0_G256_inv0 = (r00_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign z5793_assgn5793 = r10_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign m1_comar2_G4_mul5_G16_inv0_G256_inv0 = (d1_G4_mul5_G16_inv0_G256_inv0 ^ z1875_assgn1875);
    assign m2_comar2_G4_mul5_G16_inv0_G256_inv0 = (d0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign z5799_assgn5799 = r00_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign m3_comar2_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 ^ z1879_assgn1879);
    assign z5803_assgn5803 = m0_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign p2_comar2_G4_mul5_G16_inv0_G256_inv0 = (z1882_assgn1882 & m1_comar2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5807_assgn5807 = m2_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign p3_comar2_G4_mul5_G16_inv0_G256_inv0 = (m3_comar2_G4_mul5_G16_inv0_G256_inv0_reg & z1883_assgn1883);
    assign p1_comar2_G4_mul5_G16_inv0_G256_inv0 = (m0_comar2_G4_mul5_G16_inv0_G256_inv0_reg & m2_comar2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5813_assgn5813 = m1_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign p4_comar2_G4_mul5_G16_inv0_G256_inv0 = (m3_comar2_G4_mul5_G16_inv0_G256_inv0_reg & z1887_assgn1887);
    assign i0_comar2_G4_mul5_G16_inv0_G256_inv0 = (p1_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5819_assgn5819 = r1_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign i1_comar2_G4_mul5_G16_inv0_G256_inv0 = (p2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ z1891_assgn1891);
    assign z5823_assgn5823 = r2_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign i2_comar2_G4_mul5_G16_inv0_G256_inv0 = (p3_comar2_G4_mul5_G16_inv0_G256_inv0 ^ z1893_assgn1893);
    assign z5827_assgn5827 = r3_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign i3_comar2_G4_mul5_G16_inv0_G256_inv0 = (p4_comar2_G4_mul5_G16_inv0_G256_inv0 ^ z1895_assgn1895);
    assign z5831_assgn5831 = i1_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0 = (z1898_assgn1898 ^ i2_comar2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign z5835_assgn5835 = i0_comar2_G4_mul5_G16_inv0_G256_inv0;
    assign i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0 = (z1900_assgn1900 ^ i3_comar2_G4_mul5_G16_inv0_G256_inv0_reg);
    assign y1_1_comar2_G4_mul5_G16_inv0_G256_inv0 = (r00_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << dec_1_inp);
    assign z5857_assgn5857 = dec_1_inp;
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << z1919_assgn1919);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << dec_2_inp);
    assign z5867_assgn5867 = dec_2_inp;
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << z1927_assgn1927);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign r00_G16_mul1_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul1_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul1_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul1_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul1_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul1_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign z5889_assgn5889 = dec_12_inp;
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1947_assgn1947);
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign z5895_assgn5895 = dec_2_inp;
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> z1951_assgn1951);
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign z5901_assgn5901 = dec_3_inp;
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & z1955_assgn1955);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign z5939_assgn5939 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1991_assgn1991);
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign z5945_assgn5945 = dec_1_inp;
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> z1995_assgn1995);
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign z5951_assgn5951 = dec_1_inp;
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & z1999_assgn1999);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ d1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign z5993_assgn5993 = r00_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign m3_comar0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 ^ z2039_assgn2039);
    assign p2_comar0_G4_mul0_G16_mul1_G256_inv0 = (m0_comar0_G4_mul0_G16_mul1_G256_inv0_reg & m1_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z5999_assgn5999 = m2_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign p3_comar0_G4_mul0_G16_mul1_G256_inv0 = (m3_comar0_G4_mul0_G16_mul1_G256_inv0_reg & z2043_assgn2043);
    assign p1_comar0_G4_mul0_G16_mul1_G256_inv0 = (m0_comar0_G4_mul0_G16_mul1_G256_inv0_reg & m2_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6005_assgn6005 = m1_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign p4_comar0_G4_mul0_G16_mul1_G256_inv0 = (m3_comar0_G4_mul0_G16_mul1_G256_inv0_reg & z2047_assgn2047);
    assign i0_comar0_G4_mul0_G16_mul1_G256_inv0 = (p1_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign i1_comar0_G4_mul0_G16_mul1_G256_inv0 = (p2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6013_assgn6013 = r2_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign i2_comar0_G4_mul0_G16_mul1_G256_inv0 = (p3_comar0_G4_mul0_G16_mul1_G256_inv0 ^ z2053_assgn2053);
    assign z6017_assgn6017 = r3_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign i3_comar0_G4_mul0_G16_mul1_G256_inv0 = (p4_comar0_G4_mul0_G16_mul1_G256_inv0 ^ z2055_assgn2055);
    assign z6021_assgn6021 = i1_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0 = (z2058_assgn2058 ^ i2_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6025_assgn6025 = i0_comar0_G4_mul0_G16_mul1_G256_inv0;
    assign i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0 = (z2060_assgn2060 ^ i3_comar0_G4_mul0_G16_mul1_G256_inv0_reg);
    assign y1_1_comar0_G4_mul0_G16_mul1_G256_inv0 = (r00_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign z6059_assgn6059 = r00_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign m3_comar1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ z2091_assgn2091);
    assign p2_comar1_G4_mul0_G16_mul1_G256_inv0 = (m0_comar1_G4_mul0_G16_mul1_G256_inv0_reg & m1_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6065_assgn6065 = m2_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign p3_comar1_G4_mul0_G16_mul1_G256_inv0 = (m3_comar1_G4_mul0_G16_mul1_G256_inv0_reg & z2095_assgn2095);
    assign p1_comar1_G4_mul0_G16_mul1_G256_inv0 = (m0_comar1_G4_mul0_G16_mul1_G256_inv0_reg & m2_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6071_assgn6071 = m1_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign p4_comar1_G4_mul0_G16_mul1_G256_inv0 = (m3_comar1_G4_mul0_G16_mul1_G256_inv0_reg & z2099_assgn2099);
    assign i0_comar1_G4_mul0_G16_mul1_G256_inv0 = (p1_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign i1_comar1_G4_mul0_G16_mul1_G256_inv0 = (p2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6079_assgn6079 = r2_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign i2_comar1_G4_mul0_G16_mul1_G256_inv0 = (p3_comar1_G4_mul0_G16_mul1_G256_inv0 ^ z2105_assgn2105);
    assign z6083_assgn6083 = r3_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign i3_comar1_G4_mul0_G16_mul1_G256_inv0 = (p4_comar1_G4_mul0_G16_mul1_G256_inv0 ^ z2107_assgn2107);
    assign z6087_assgn6087 = i1_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0 = (z2110_assgn2110 ^ i2_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6091_assgn6091 = i0_comar1_G4_mul0_G16_mul1_G256_inv0;
    assign i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0 = (z2112_assgn2112 ^ i3_comar1_G4_mul0_G16_mul1_G256_inv0_reg);
    assign y1_1_comar1_G4_mul0_G16_mul1_G256_inv0 = (r00_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul1_G256_inv0 = (d1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul1_G256_inv0 = (d0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign z6129_assgn6129 = r00_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign m3_comar2_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 ^ z2147_assgn2147);
    assign p2_comar2_G4_mul0_G16_mul1_G256_inv0 = (m0_comar2_G4_mul0_G16_mul1_G256_inv0_reg & m1_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6135_assgn6135 = m2_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign p3_comar2_G4_mul0_G16_mul1_G256_inv0 = (m3_comar2_G4_mul0_G16_mul1_G256_inv0_reg & z2151_assgn2151);
    assign p1_comar2_G4_mul0_G16_mul1_G256_inv0 = (m0_comar2_G4_mul0_G16_mul1_G256_inv0_reg & m2_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6141_assgn6141 = m1_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign p4_comar2_G4_mul0_G16_mul1_G256_inv0 = (m3_comar2_G4_mul0_G16_mul1_G256_inv0_reg & z2155_assgn2155);
    assign i0_comar2_G4_mul0_G16_mul1_G256_inv0 = (p1_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign i1_comar2_G4_mul0_G16_mul1_G256_inv0 = (p2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6149_assgn6149 = r2_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign i2_comar2_G4_mul0_G16_mul1_G256_inv0 = (p3_comar2_G4_mul0_G16_mul1_G256_inv0 ^ z2161_assgn2161);
    assign z6153_assgn6153 = r3_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign i3_comar2_G4_mul0_G16_mul1_G256_inv0 = (p4_comar2_G4_mul0_G16_mul1_G256_inv0 ^ z2163_assgn2163);
    assign z6157_assgn6157 = i1_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0 = (z2166_assgn2166 ^ i2_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign z6161_assgn6161 = i0_comar2_G4_mul0_G16_mul1_G256_inv0;
    assign i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0 = (z2168_assgn2168 ^ i3_comar2_G4_mul0_G16_mul1_G256_inv0_reg);
    assign y1_1_comar2_G4_mul0_G16_mul1_G256_inv0 = (r00_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << dec_1_inp);
    assign z6183_assgn6183 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << z2187_assgn2187);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_2_inp);
    assign z6193_assgn6193 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z2195_assgn2195);
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign z6199_assgn6199 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> z2199_assgn2199);
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_1_inp);
    assign z6205_assgn6205 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & z2203_assgn2203);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign z6217_assgn6217 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << z2213_assgn2213);
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << dec_1_inp);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_2_inp);
    assign z6241_assgn6241 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z2235_assgn2235);
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign z6247_assgn6247 = dec_1_inp;
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> z2239_assgn2239);
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_1_inp);
    assign z6253_assgn6253 = dec_1_inp;
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & z2243_assgn2243);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ d1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul1_G256_inv0 = (cxord_1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul1_G256_inv0 = (cxord_0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign z6295_assgn6295 = r00_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign m3_comar0_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 ^ z2283_assgn2283);
    assign p2_comar0_G4_mul1_G16_mul1_G256_inv0 = (m0_comar0_G4_mul1_G16_mul1_G256_inv0_reg & m1_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6301_assgn6301 = m2_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign p3_comar0_G4_mul1_G16_mul1_G256_inv0 = (m3_comar0_G4_mul1_G16_mul1_G256_inv0_reg & z2287_assgn2287);
    assign p1_comar0_G4_mul1_G16_mul1_G256_inv0 = (m0_comar0_G4_mul1_G16_mul1_G256_inv0_reg & m2_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6307_assgn6307 = m1_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign p4_comar0_G4_mul1_G16_mul1_G256_inv0 = (m3_comar0_G4_mul1_G16_mul1_G256_inv0_reg & z2291_assgn2291);
    assign i0_comar0_G4_mul1_G16_mul1_G256_inv0 = (p1_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign i1_comar0_G4_mul1_G16_mul1_G256_inv0 = (p2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6315_assgn6315 = r2_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign i2_comar0_G4_mul1_G16_mul1_G256_inv0 = (p3_comar0_G4_mul1_G16_mul1_G256_inv0 ^ z2297_assgn2297);
    assign z6319_assgn6319 = r3_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign i3_comar0_G4_mul1_G16_mul1_G256_inv0 = (p4_comar0_G4_mul1_G16_mul1_G256_inv0 ^ z2299_assgn2299);
    assign z6323_assgn6323 = i1_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0 = (z2302_assgn2302 ^ i2_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6327_assgn6327 = i0_comar0_G4_mul1_G16_mul1_G256_inv0;
    assign i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0 = (z2304_assgn2304 ^ i3_comar0_G4_mul1_G16_mul1_G256_inv0_reg);
    assign y1_1_comar0_G4_mul1_G16_mul1_G256_inv0 = (r00_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign z6361_assgn6361 = r00_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign m3_comar1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ z2335_assgn2335);
    assign p2_comar1_G4_mul1_G16_mul1_G256_inv0 = (m0_comar1_G4_mul1_G16_mul1_G256_inv0_reg & m1_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6367_assgn6367 = m2_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign p3_comar1_G4_mul1_G16_mul1_G256_inv0 = (m3_comar1_G4_mul1_G16_mul1_G256_inv0_reg & z2339_assgn2339);
    assign p1_comar1_G4_mul1_G16_mul1_G256_inv0 = (m0_comar1_G4_mul1_G16_mul1_G256_inv0_reg & m2_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6373_assgn6373 = m1_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign p4_comar1_G4_mul1_G16_mul1_G256_inv0 = (m3_comar1_G4_mul1_G16_mul1_G256_inv0_reg & z2343_assgn2343);
    assign i0_comar1_G4_mul1_G16_mul1_G256_inv0 = (p1_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign i1_comar1_G4_mul1_G16_mul1_G256_inv0 = (p2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6381_assgn6381 = r2_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign i2_comar1_G4_mul1_G16_mul1_G256_inv0 = (p3_comar1_G4_mul1_G16_mul1_G256_inv0 ^ z2349_assgn2349);
    assign z6385_assgn6385 = r3_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign i3_comar1_G4_mul1_G16_mul1_G256_inv0 = (p4_comar1_G4_mul1_G16_mul1_G256_inv0 ^ z2351_assgn2351);
    assign z6389_assgn6389 = i1_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0 = (z2354_assgn2354 ^ i2_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6393_assgn6393 = i0_comar1_G4_mul1_G16_mul1_G256_inv0;
    assign i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0 = (z2356_assgn2356 ^ i3_comar1_G4_mul1_G16_mul1_G256_inv0_reg);
    assign y1_1_comar1_G4_mul1_G16_mul1_G256_inv0 = (r00_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul1_G256_inv0 = (d1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul1_G256_inv0 = (d0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign z6431_assgn6431 = r00_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign m3_comar2_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 ^ z2391_assgn2391);
    assign p2_comar2_G4_mul1_G16_mul1_G256_inv0 = (m0_comar2_G4_mul1_G16_mul1_G256_inv0_reg & m1_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6437_assgn6437 = m2_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign p3_comar2_G4_mul1_G16_mul1_G256_inv0 = (m3_comar2_G4_mul1_G16_mul1_G256_inv0_reg & z2395_assgn2395);
    assign p1_comar2_G4_mul1_G16_mul1_G256_inv0 = (m0_comar2_G4_mul1_G16_mul1_G256_inv0_reg & m2_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6443_assgn6443 = m1_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign p4_comar2_G4_mul1_G16_mul1_G256_inv0 = (m3_comar2_G4_mul1_G16_mul1_G256_inv0_reg & z2399_assgn2399);
    assign i0_comar2_G4_mul1_G16_mul1_G256_inv0 = (p1_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign i1_comar2_G4_mul1_G16_mul1_G256_inv0 = (p2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6451_assgn6451 = r2_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign i2_comar2_G4_mul1_G16_mul1_G256_inv0 = (p3_comar2_G4_mul1_G16_mul1_G256_inv0 ^ z2405_assgn2405);
    assign z6455_assgn6455 = r3_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign i3_comar2_G4_mul1_G16_mul1_G256_inv0 = (p4_comar2_G4_mul1_G16_mul1_G256_inv0 ^ z2407_assgn2407);
    assign z6459_assgn6459 = i1_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0 = (z2410_assgn2410 ^ i2_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign z6463_assgn6463 = i0_comar2_G4_mul1_G16_mul1_G256_inv0;
    assign i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0 = (z2412_assgn2412 ^ i3_comar2_G4_mul1_G16_mul1_G256_inv0_reg);
    assign y1_1_comar2_G4_mul1_G16_mul1_G256_inv0 = (r00_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << dec_1_inp);
    assign z6485_assgn6485 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << z2431_assgn2431);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_2_inp);
    assign z6511_assgn6511 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z2455_assgn2455);
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign z6517_assgn6517 = dec_1_inp;
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> z2459_assgn2459);
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_1_inp);
    assign z6523_assgn6523 = dec_1_inp;
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & z2463_assgn2463);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ d1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul1_G256_inv0 = (cxord_1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul1_G256_inv0 = (cxord_0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign z6565_assgn6565 = r00_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign m3_comar0_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 ^ z2503_assgn2503);
    assign p2_comar0_G4_mul2_G16_mul1_G256_inv0 = (m0_comar0_G4_mul2_G16_mul1_G256_inv0_reg & m1_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6571_assgn6571 = m2_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign p3_comar0_G4_mul2_G16_mul1_G256_inv0 = (m3_comar0_G4_mul2_G16_mul1_G256_inv0_reg & z2507_assgn2507);
    assign p1_comar0_G4_mul2_G16_mul1_G256_inv0 = (m0_comar0_G4_mul2_G16_mul1_G256_inv0_reg & m2_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6577_assgn6577 = m1_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign p4_comar0_G4_mul2_G16_mul1_G256_inv0 = (m3_comar0_G4_mul2_G16_mul1_G256_inv0_reg & z2511_assgn2511);
    assign i0_comar0_G4_mul2_G16_mul1_G256_inv0 = (p1_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign i1_comar0_G4_mul2_G16_mul1_G256_inv0 = (p2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6585_assgn6585 = r2_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign i2_comar0_G4_mul2_G16_mul1_G256_inv0 = (p3_comar0_G4_mul2_G16_mul1_G256_inv0 ^ z2517_assgn2517);
    assign z6589_assgn6589 = r3_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign i3_comar0_G4_mul2_G16_mul1_G256_inv0 = (p4_comar0_G4_mul2_G16_mul1_G256_inv0 ^ z2519_assgn2519);
    assign z6593_assgn6593 = i1_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0 = (z2522_assgn2522 ^ i2_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6597_assgn6597 = i0_comar0_G4_mul2_G16_mul1_G256_inv0;
    assign i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0 = (z2524_assgn2524 ^ i3_comar0_G4_mul2_G16_mul1_G256_inv0_reg);
    assign y1_1_comar0_G4_mul2_G16_mul1_G256_inv0 = (r00_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign z6631_assgn6631 = r00_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign m3_comar1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ z2555_assgn2555);
    assign p2_comar1_G4_mul2_G16_mul1_G256_inv0 = (m0_comar1_G4_mul2_G16_mul1_G256_inv0_reg & m1_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6637_assgn6637 = m2_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign p3_comar1_G4_mul2_G16_mul1_G256_inv0 = (m3_comar1_G4_mul2_G16_mul1_G256_inv0_reg & z2559_assgn2559);
    assign p1_comar1_G4_mul2_G16_mul1_G256_inv0 = (m0_comar1_G4_mul2_G16_mul1_G256_inv0_reg & m2_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6643_assgn6643 = m1_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign p4_comar1_G4_mul2_G16_mul1_G256_inv0 = (m3_comar1_G4_mul2_G16_mul1_G256_inv0_reg & z2563_assgn2563);
    assign i0_comar1_G4_mul2_G16_mul1_G256_inv0 = (p1_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign i1_comar1_G4_mul2_G16_mul1_G256_inv0 = (p2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6651_assgn6651 = r2_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign i2_comar1_G4_mul2_G16_mul1_G256_inv0 = (p3_comar1_G4_mul2_G16_mul1_G256_inv0 ^ z2569_assgn2569);
    assign z6655_assgn6655 = r3_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign i3_comar1_G4_mul2_G16_mul1_G256_inv0 = (p4_comar1_G4_mul2_G16_mul1_G256_inv0 ^ z2571_assgn2571);
    assign z6659_assgn6659 = i1_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0 = (z2574_assgn2574 ^ i2_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6663_assgn6663 = i0_comar1_G4_mul2_G16_mul1_G256_inv0;
    assign i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0 = (z2576_assgn2576 ^ i3_comar1_G4_mul2_G16_mul1_G256_inv0_reg);
    assign y1_1_comar1_G4_mul2_G16_mul1_G256_inv0 = (r00_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul1_G256_inv0 = (d1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul1_G256_inv0 = (d0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign z6701_assgn6701 = r00_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign m3_comar2_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 ^ z2611_assgn2611);
    assign p2_comar2_G4_mul2_G16_mul1_G256_inv0 = (m0_comar2_G4_mul2_G16_mul1_G256_inv0_reg & m1_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6707_assgn6707 = m2_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign p3_comar2_G4_mul2_G16_mul1_G256_inv0 = (m3_comar2_G4_mul2_G16_mul1_G256_inv0_reg & z2615_assgn2615);
    assign p1_comar2_G4_mul2_G16_mul1_G256_inv0 = (m0_comar2_G4_mul2_G16_mul1_G256_inv0_reg & m2_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6713_assgn6713 = m1_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign p4_comar2_G4_mul2_G16_mul1_G256_inv0 = (m3_comar2_G4_mul2_G16_mul1_G256_inv0_reg & z2619_assgn2619);
    assign i0_comar2_G4_mul2_G16_mul1_G256_inv0 = (p1_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign i1_comar2_G4_mul2_G16_mul1_G256_inv0 = (p2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6721_assgn6721 = r2_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign i2_comar2_G4_mul2_G16_mul1_G256_inv0 = (p3_comar2_G4_mul2_G16_mul1_G256_inv0 ^ z2625_assgn2625);
    assign z6725_assgn6725 = r3_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign i3_comar2_G4_mul2_G16_mul1_G256_inv0 = (p4_comar2_G4_mul2_G16_mul1_G256_inv0 ^ z2627_assgn2627);
    assign z6729_assgn6729 = i1_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0 = (z2630_assgn2630 ^ i2_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign z6733_assgn6733 = i0_comar2_G4_mul2_G16_mul1_G256_inv0;
    assign i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0 = (z2632_assgn2632 ^ i3_comar2_G4_mul2_G16_mul1_G256_inv0_reg);
    assign y1_1_comar2_G4_mul2_G16_mul1_G256_inv0 = (r00_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << dec_1_inp);
    assign z6755_assgn6755 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << z2651_assgn2651);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << dec_2_inp);
    assign z6769_assgn6769 = dec_2_inp;
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << z2663_assgn2663);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign r00_G16_mul2_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul2_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul2_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul2_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul2_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul2_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign z6791_assgn6791 = dec_12_inp;
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2683_assgn2683);
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign z6797_assgn6797 = dec_2_inp;
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> z2687_assgn2687);
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign z6803_assgn6803 = dec_3_inp;
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & z2691_assgn2691);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign z6841_assgn6841 = dec_2_inp;
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2727_assgn2727);
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign z6847_assgn6847 = dec_1_inp;
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> z2731_assgn2731);
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign z6853_assgn6853 = dec_1_inp;
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & z2735_assgn2735);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ d1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign z6895_assgn6895 = r00_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign m3_comar0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 ^ z2775_assgn2775);
    assign p2_comar0_G4_mul0_G16_mul2_G256_inv0 = (m0_comar0_G4_mul0_G16_mul2_G256_inv0_reg & m1_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6901_assgn6901 = m2_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign p3_comar0_G4_mul0_G16_mul2_G256_inv0 = (m3_comar0_G4_mul0_G16_mul2_G256_inv0_reg & z2779_assgn2779);
    assign p1_comar0_G4_mul0_G16_mul2_G256_inv0 = (m0_comar0_G4_mul0_G16_mul2_G256_inv0_reg & m2_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6907_assgn6907 = m1_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign p4_comar0_G4_mul0_G16_mul2_G256_inv0 = (m3_comar0_G4_mul0_G16_mul2_G256_inv0_reg & z2783_assgn2783);
    assign i0_comar0_G4_mul0_G16_mul2_G256_inv0 = (p1_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign i1_comar0_G4_mul0_G16_mul2_G256_inv0 = (p2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6915_assgn6915 = r2_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign i2_comar0_G4_mul0_G16_mul2_G256_inv0 = (p3_comar0_G4_mul0_G16_mul2_G256_inv0 ^ z2789_assgn2789);
    assign z6919_assgn6919 = r3_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign i3_comar0_G4_mul0_G16_mul2_G256_inv0 = (p4_comar0_G4_mul0_G16_mul2_G256_inv0 ^ z2791_assgn2791);
    assign z6923_assgn6923 = i1_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0 = (z2794_assgn2794 ^ i2_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6927_assgn6927 = i0_comar0_G4_mul0_G16_mul2_G256_inv0;
    assign i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0 = (z2796_assgn2796 ^ i3_comar0_G4_mul0_G16_mul2_G256_inv0_reg);
    assign y1_1_comar0_G4_mul0_G16_mul2_G256_inv0 = (r00_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign z6961_assgn6961 = r00_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign m3_comar1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ z2827_assgn2827);
    assign p2_comar1_G4_mul0_G16_mul2_G256_inv0 = (m0_comar1_G4_mul0_G16_mul2_G256_inv0_reg & m1_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6967_assgn6967 = m2_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign p3_comar1_G4_mul0_G16_mul2_G256_inv0 = (m3_comar1_G4_mul0_G16_mul2_G256_inv0_reg & z2831_assgn2831);
    assign p1_comar1_G4_mul0_G16_mul2_G256_inv0 = (m0_comar1_G4_mul0_G16_mul2_G256_inv0_reg & m2_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6973_assgn6973 = m1_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign p4_comar1_G4_mul0_G16_mul2_G256_inv0 = (m3_comar1_G4_mul0_G16_mul2_G256_inv0_reg & z2835_assgn2835);
    assign i0_comar1_G4_mul0_G16_mul2_G256_inv0 = (p1_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign i1_comar1_G4_mul0_G16_mul2_G256_inv0 = (p2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6981_assgn6981 = r2_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign i2_comar1_G4_mul0_G16_mul2_G256_inv0 = (p3_comar1_G4_mul0_G16_mul2_G256_inv0 ^ z2841_assgn2841);
    assign z6985_assgn6985 = r3_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign i3_comar1_G4_mul0_G16_mul2_G256_inv0 = (p4_comar1_G4_mul0_G16_mul2_G256_inv0 ^ z2843_assgn2843);
    assign z6989_assgn6989 = i1_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0 = (z2846_assgn2846 ^ i2_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z6993_assgn6993 = i0_comar1_G4_mul0_G16_mul2_G256_inv0;
    assign i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0 = (z2848_assgn2848 ^ i3_comar1_G4_mul0_G16_mul2_G256_inv0_reg);
    assign y1_1_comar1_G4_mul0_G16_mul2_G256_inv0 = (r00_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul2_G256_inv0 = (d1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul2_G256_inv0 = (d0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign z7031_assgn7031 = r00_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign m3_comar2_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 ^ z2883_assgn2883);
    assign p2_comar2_G4_mul0_G16_mul2_G256_inv0 = (m0_comar2_G4_mul0_G16_mul2_G256_inv0_reg & m1_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z7037_assgn7037 = m2_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign p3_comar2_G4_mul0_G16_mul2_G256_inv0 = (m3_comar2_G4_mul0_G16_mul2_G256_inv0_reg & z2887_assgn2887);
    assign p1_comar2_G4_mul0_G16_mul2_G256_inv0 = (m0_comar2_G4_mul0_G16_mul2_G256_inv0_reg & m2_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z7043_assgn7043 = m1_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign p4_comar2_G4_mul0_G16_mul2_G256_inv0 = (m3_comar2_G4_mul0_G16_mul2_G256_inv0_reg & z2891_assgn2891);
    assign i0_comar2_G4_mul0_G16_mul2_G256_inv0 = (p1_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign i1_comar2_G4_mul0_G16_mul2_G256_inv0 = (p2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z7051_assgn7051 = r2_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign i2_comar2_G4_mul0_G16_mul2_G256_inv0 = (p3_comar2_G4_mul0_G16_mul2_G256_inv0 ^ z2897_assgn2897);
    assign z7055_assgn7055 = r3_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign i3_comar2_G4_mul0_G16_mul2_G256_inv0 = (p4_comar2_G4_mul0_G16_mul2_G256_inv0 ^ z2899_assgn2899);
    assign z7059_assgn7059 = i1_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0 = (z2902_assgn2902 ^ i2_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign z7063_assgn7063 = i0_comar2_G4_mul0_G16_mul2_G256_inv0;
    assign i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0 = (z2904_assgn2904 ^ i3_comar2_G4_mul0_G16_mul2_G256_inv0_reg);
    assign y1_1_comar2_G4_mul0_G16_mul2_G256_inv0 = (r00_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << dec_1_inp);
    assign z7085_assgn7085 = dec_1_inp;
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << z2923_assgn2923);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_2_inp);
    assign z7095_assgn7095 = dec_2_inp;
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2931_assgn2931);
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign z7101_assgn7101 = dec_1_inp;
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> z2935_assgn2935);
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_1_inp);
    assign z7107_assgn7107 = dec_1_inp;
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & z2939_assgn2939);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign z7119_assgn7119 = dec_1_inp;
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << z2949_assgn2949);
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << dec_1_inp);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_2_inp);
    assign z7143_assgn7143 = dec_2_inp;
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2971_assgn2971);
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign z7149_assgn7149 = dec_1_inp;
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> z2975_assgn2975);
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_1_inp);
    assign z7155_assgn7155 = dec_1_inp;
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & z2979_assgn2979);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ d1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul2_G256_inv0 = (cxord_1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul2_G256_inv0 = (cxord_0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign z7197_assgn7197 = r00_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign m3_comar0_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 ^ z3019_assgn3019);
    assign p2_comar0_G4_mul1_G16_mul2_G256_inv0 = (m0_comar0_G4_mul1_G16_mul2_G256_inv0_reg & m1_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7203_assgn7203 = m2_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign p3_comar0_G4_mul1_G16_mul2_G256_inv0 = (m3_comar0_G4_mul1_G16_mul2_G256_inv0_reg & z3023_assgn3023);
    assign p1_comar0_G4_mul1_G16_mul2_G256_inv0 = (m0_comar0_G4_mul1_G16_mul2_G256_inv0_reg & m2_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7209_assgn7209 = m1_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign p4_comar0_G4_mul1_G16_mul2_G256_inv0 = (m3_comar0_G4_mul1_G16_mul2_G256_inv0_reg & z3027_assgn3027);
    assign i0_comar0_G4_mul1_G16_mul2_G256_inv0 = (p1_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign i1_comar0_G4_mul1_G16_mul2_G256_inv0 = (p2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7217_assgn7217 = r2_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign i2_comar0_G4_mul1_G16_mul2_G256_inv0 = (p3_comar0_G4_mul1_G16_mul2_G256_inv0 ^ z3033_assgn3033);
    assign z7221_assgn7221 = r3_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign i3_comar0_G4_mul1_G16_mul2_G256_inv0 = (p4_comar0_G4_mul1_G16_mul2_G256_inv0 ^ z3035_assgn3035);
    assign z7225_assgn7225 = i1_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0 = (z3038_assgn3038 ^ i2_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7229_assgn7229 = i0_comar0_G4_mul1_G16_mul2_G256_inv0;
    assign i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0 = (z3040_assgn3040 ^ i3_comar0_G4_mul1_G16_mul2_G256_inv0_reg);
    assign y1_1_comar0_G4_mul1_G16_mul2_G256_inv0 = (r00_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign z7263_assgn7263 = r00_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign m3_comar1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ z3071_assgn3071);
    assign p2_comar1_G4_mul1_G16_mul2_G256_inv0 = (m0_comar1_G4_mul1_G16_mul2_G256_inv0_reg & m1_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7269_assgn7269 = m2_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign p3_comar1_G4_mul1_G16_mul2_G256_inv0 = (m3_comar1_G4_mul1_G16_mul2_G256_inv0_reg & z3075_assgn3075);
    assign p1_comar1_G4_mul1_G16_mul2_G256_inv0 = (m0_comar1_G4_mul1_G16_mul2_G256_inv0_reg & m2_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7275_assgn7275 = m1_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign p4_comar1_G4_mul1_G16_mul2_G256_inv0 = (m3_comar1_G4_mul1_G16_mul2_G256_inv0_reg & z3079_assgn3079);
    assign i0_comar1_G4_mul1_G16_mul2_G256_inv0 = (p1_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign i1_comar1_G4_mul1_G16_mul2_G256_inv0 = (p2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7283_assgn7283 = r2_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign i2_comar1_G4_mul1_G16_mul2_G256_inv0 = (p3_comar1_G4_mul1_G16_mul2_G256_inv0 ^ z3085_assgn3085);
    assign z7287_assgn7287 = r3_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign i3_comar1_G4_mul1_G16_mul2_G256_inv0 = (p4_comar1_G4_mul1_G16_mul2_G256_inv0 ^ z3087_assgn3087);
    assign z7291_assgn7291 = i1_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0 = (z3090_assgn3090 ^ i2_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7295_assgn7295 = i0_comar1_G4_mul1_G16_mul2_G256_inv0;
    assign i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0 = (z3092_assgn3092 ^ i3_comar1_G4_mul1_G16_mul2_G256_inv0_reg);
    assign y1_1_comar1_G4_mul1_G16_mul2_G256_inv0 = (r00_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul2_G256_inv0 = (d1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul2_G256_inv0 = (d0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign z7333_assgn7333 = r00_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign m3_comar2_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 ^ z3127_assgn3127);
    assign p2_comar2_G4_mul1_G16_mul2_G256_inv0 = (m0_comar2_G4_mul1_G16_mul2_G256_inv0_reg & m1_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7339_assgn7339 = m2_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign p3_comar2_G4_mul1_G16_mul2_G256_inv0 = (m3_comar2_G4_mul1_G16_mul2_G256_inv0_reg & z3131_assgn3131);
    assign p1_comar2_G4_mul1_G16_mul2_G256_inv0 = (m0_comar2_G4_mul1_G16_mul2_G256_inv0_reg & m2_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7345_assgn7345 = m1_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign p4_comar2_G4_mul1_G16_mul2_G256_inv0 = (m3_comar2_G4_mul1_G16_mul2_G256_inv0_reg & z3135_assgn3135);
    assign i0_comar2_G4_mul1_G16_mul2_G256_inv0 = (p1_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign i1_comar2_G4_mul1_G16_mul2_G256_inv0 = (p2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7353_assgn7353 = r2_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign i2_comar2_G4_mul1_G16_mul2_G256_inv0 = (p3_comar2_G4_mul1_G16_mul2_G256_inv0 ^ z3141_assgn3141);
    assign z7357_assgn7357 = r3_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign i3_comar2_G4_mul1_G16_mul2_G256_inv0 = (p4_comar2_G4_mul1_G16_mul2_G256_inv0 ^ z3143_assgn3143);
    assign z7361_assgn7361 = i1_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0 = (z3146_assgn3146 ^ i2_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign z7365_assgn7365 = i0_comar2_G4_mul1_G16_mul2_G256_inv0;
    assign i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0 = (z3148_assgn3148 ^ i3_comar2_G4_mul1_G16_mul2_G256_inv0_reg);
    assign y1_1_comar2_G4_mul1_G16_mul2_G256_inv0 = (r00_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << dec_1_inp);
    assign z7387_assgn7387 = dec_1_inp;
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << z3167_assgn3167);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_2_inp);
    assign z7413_assgn7413 = dec_2_inp;
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z3191_assgn3191);
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign z7419_assgn7419 = dec_1_inp;
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> z3195_assgn3195);
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_1_inp);
    assign z7425_assgn7425 = dec_1_inp;
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & z3199_assgn3199);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ d1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul2_G256_inv0 = (cxord_1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul2_G256_inv0 = (cxord_0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign z7467_assgn7467 = r00_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign m3_comar0_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 ^ z3239_assgn3239);
    assign p2_comar0_G4_mul2_G16_mul2_G256_inv0 = (m0_comar0_G4_mul2_G16_mul2_G256_inv0_reg & m1_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7473_assgn7473 = m2_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign p3_comar0_G4_mul2_G16_mul2_G256_inv0 = (m3_comar0_G4_mul2_G16_mul2_G256_inv0_reg & z3243_assgn3243);
    assign p1_comar0_G4_mul2_G16_mul2_G256_inv0 = (m0_comar0_G4_mul2_G16_mul2_G256_inv0_reg & m2_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7479_assgn7479 = m1_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign p4_comar0_G4_mul2_G16_mul2_G256_inv0 = (m3_comar0_G4_mul2_G16_mul2_G256_inv0_reg & z3247_assgn3247);
    assign i0_comar0_G4_mul2_G16_mul2_G256_inv0 = (p1_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign i1_comar0_G4_mul2_G16_mul2_G256_inv0 = (p2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7487_assgn7487 = r2_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign i2_comar0_G4_mul2_G16_mul2_G256_inv0 = (p3_comar0_G4_mul2_G16_mul2_G256_inv0 ^ z3253_assgn3253);
    assign z7491_assgn7491 = r3_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign i3_comar0_G4_mul2_G16_mul2_G256_inv0 = (p4_comar0_G4_mul2_G16_mul2_G256_inv0 ^ z3255_assgn3255);
    assign z7495_assgn7495 = i1_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0 = (z3258_assgn3258 ^ i2_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7499_assgn7499 = i0_comar0_G4_mul2_G16_mul2_G256_inv0;
    assign i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0 = (z3260_assgn3260 ^ i3_comar0_G4_mul2_G16_mul2_G256_inv0_reg);
    assign y1_1_comar0_G4_mul2_G16_mul2_G256_inv0 = (r00_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign z7533_assgn7533 = r00_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign m3_comar1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ z3291_assgn3291);
    assign p2_comar1_G4_mul2_G16_mul2_G256_inv0 = (m0_comar1_G4_mul2_G16_mul2_G256_inv0_reg & m1_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7539_assgn7539 = m2_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign p3_comar1_G4_mul2_G16_mul2_G256_inv0 = (m3_comar1_G4_mul2_G16_mul2_G256_inv0_reg & z3295_assgn3295);
    assign p1_comar1_G4_mul2_G16_mul2_G256_inv0 = (m0_comar1_G4_mul2_G16_mul2_G256_inv0_reg & m2_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7545_assgn7545 = m1_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign p4_comar1_G4_mul2_G16_mul2_G256_inv0 = (m3_comar1_G4_mul2_G16_mul2_G256_inv0_reg & z3299_assgn3299);
    assign i0_comar1_G4_mul2_G16_mul2_G256_inv0 = (p1_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign i1_comar1_G4_mul2_G16_mul2_G256_inv0 = (p2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7553_assgn7553 = r2_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign i2_comar1_G4_mul2_G16_mul2_G256_inv0 = (p3_comar1_G4_mul2_G16_mul2_G256_inv0 ^ z3305_assgn3305);
    assign z7557_assgn7557 = r3_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign i3_comar1_G4_mul2_G16_mul2_G256_inv0 = (p4_comar1_G4_mul2_G16_mul2_G256_inv0 ^ z3307_assgn3307);
    assign z7561_assgn7561 = i1_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0 = (z3310_assgn3310 ^ i2_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7565_assgn7565 = i0_comar1_G4_mul2_G16_mul2_G256_inv0;
    assign i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0 = (z3312_assgn3312 ^ i3_comar1_G4_mul2_G16_mul2_G256_inv0_reg);
    assign y1_1_comar1_G4_mul2_G16_mul2_G256_inv0 = (r00_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul2_G256_inv0 = (d1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul2_G256_inv0 = (d0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign z7603_assgn7603 = r00_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign m3_comar2_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 ^ z3347_assgn3347);
    assign p2_comar2_G4_mul2_G16_mul2_G256_inv0 = (m0_comar2_G4_mul2_G16_mul2_G256_inv0_reg & m1_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7609_assgn7609 = m2_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign p3_comar2_G4_mul2_G16_mul2_G256_inv0 = (m3_comar2_G4_mul2_G16_mul2_G256_inv0_reg & z3351_assgn3351);
    assign p1_comar2_G4_mul2_G16_mul2_G256_inv0 = (m0_comar2_G4_mul2_G16_mul2_G256_inv0_reg & m2_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7615_assgn7615 = m1_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign p4_comar2_G4_mul2_G16_mul2_G256_inv0 = (m3_comar2_G4_mul2_G16_mul2_G256_inv0_reg & z3355_assgn3355);
    assign i0_comar2_G4_mul2_G16_mul2_G256_inv0 = (p1_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign i1_comar2_G4_mul2_G16_mul2_G256_inv0 = (p2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7623_assgn7623 = r2_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign i2_comar2_G4_mul2_G16_mul2_G256_inv0 = (p3_comar2_G4_mul2_G16_mul2_G256_inv0 ^ z3361_assgn3361);
    assign z7627_assgn7627 = r3_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign i3_comar2_G4_mul2_G16_mul2_G256_inv0 = (p4_comar2_G4_mul2_G16_mul2_G256_inv0 ^ z3363_assgn3363);
    assign z7631_assgn7631 = i1_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0 = (z3366_assgn3366 ^ i2_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign z7635_assgn7635 = i0_comar2_G4_mul2_G16_mul2_G256_inv0;
    assign i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0 = (z3368_assgn3368 ^ i3_comar2_G4_mul2_G16_mul2_G256_inv0_reg);
    assign y1_1_comar2_G4_mul2_G16_mul2_G256_inv0 = (r00_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << dec_1_inp);
    assign z7657_assgn7657 = dec_1_inp;
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << z3387_assgn3387);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << dec_2_inp);
    assign z7671_assgn7671 = dec_2_inp;
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << z3399_assgn3399);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << dec_4_inp);
    assign z7681_assgn7681 = dec_4_inp;
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << z3407_assgn3407);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign cond1_G256_newbasis1 = (t4 & dec_1_inp);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * yxorb1_G256_newbasis1);
    assign tempyIntoNegCond1_G256_newbasis1 = (tempy1_G256_newbasis1 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempyIntoNegCond1_G256_newbasis1);
    assign x1_G256_newbasis1 = (t4 >> dec_1_inp);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & dec_1_inp);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ dec_3_inp);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempyIntoNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempyIntoNegCond2_G256_newbasis1);
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> dec_1_inp);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & dec_1_inp);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ dec_4_inp);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempyIntoNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempyIntoNegCond3_G256_newbasis1);
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> dec_1_inp);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & dec_1_inp);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ dec_220_inp);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempyIntoNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempyIntoNegCond4_G256_newbasis1);
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> dec_1_inp);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & dec_1_inp);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ dec_11_inp);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempyIntoNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempyIntoNegCond5_G256_newbasis1);
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> dec_1_inp);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & dec_1_inp);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ dec_158_inp);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempyIntoNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempyIntoNegCond6_G256_newbasis1);
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> dec_1_inp);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & dec_1_inp);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ dec_45_inp);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempyIntoNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempyIntoNegCond7_G256_newbasis1);
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> dec_1_inp);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & dec_1_inp);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ dec_88_inp);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempyIntoNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempyIntoNegCond8_G256_newbasis1);
    assign z7817_assgn7817 = (x7_G256_newbasis1 >> dec_1_inp);
    assign t6 = y8_G256_newbasis1;
    assign z_y_G256_newbasis1 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z7825_assgn7825 = dec_1_inp;
    assign z_cond1_G256_newbasis1 = (t5 & z3549_assgn3549);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z7833_assgn7833 = z_yxorb1_G256_newbasis1;
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z3555_assgn3555);
    assign z7837_assgn7837 = z_tempy1_G256_newbasis1;
    assign z_tempyIntoNegCond1_G256_newbasis1 = (z3558_assgn3558 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempyIntoNegCond1_G256_newbasis1);
    assign z7843_assgn7843 = dec_1_inp;
    assign z_x1_G256_newbasis1 = (t5 >> z3561_assgn3561);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z7849_assgn7849 = dec_1_inp;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & z3565_assgn3565);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z7855_assgn7855 = dec_3_inp;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ z3569_assgn3569);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempyIntoNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempyIntoNegCond2_G256_newbasis1);
    assign z7865_assgn7865 = dec_1_inp;
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> z3577_assgn3577);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z7871_assgn7871 = dec_1_inp;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & z3581_assgn3581);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z7877_assgn7877 = dec_4_inp;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ z3585_assgn3585);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempyIntoNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempyIntoNegCond3_G256_newbasis1);
    assign z7887_assgn7887 = dec_1_inp;
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> z3593_assgn3593);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z7893_assgn7893 = dec_1_inp;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & z3597_assgn3597);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z7899_assgn7899 = dec_220_inp;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ z3601_assgn3601);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempyIntoNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempyIntoNegCond4_G256_newbasis1);
    assign z7909_assgn7909 = dec_1_inp;
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> z3609_assgn3609);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z7915_assgn7915 = dec_1_inp;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & z3613_assgn3613);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z7921_assgn7921 = dec_11_inp;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ z3617_assgn3617);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempyIntoNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempyIntoNegCond5_G256_newbasis1);
    assign z7931_assgn7931 = dec_1_inp;
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> z3625_assgn3625);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z7937_assgn7937 = dec_1_inp;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & z3629_assgn3629);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z7943_assgn7943 = dec_158_inp;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ z3633_assgn3633);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempyIntoNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempyIntoNegCond6_G256_newbasis1);
    assign z7953_assgn7953 = dec_1_inp;
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> z3641_assgn3641);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z7959_assgn7959 = dec_1_inp;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & z3645_assgn3645);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z7965_assgn7965 = dec_45_inp;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ z3649_assgn3649);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempyIntoNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempyIntoNegCond7_G256_newbasis1);
    assign z7975_assgn7975 = dec_1_inp;
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> z3657_assgn3657);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z7981_assgn7981 = dec_1_inp;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & z3661_assgn3661);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z7987_assgn7987 = dec_88_inp;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ z3665_assgn3665);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempyIntoNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempyIntoNegCond8_G256_newbasis1);
    assign z7997_assgn7997 = dec_1_inp;
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> z3673_assgn3673);
    assign t7 = z_y8_G256_newbasis1;
    assign z8003_assgn8003 = (t6 ^ dec_99_inp);

    always @(posedge clk) begin
        z3873_assgn38730 <= z3873_assgn3873;
        z3873_assgn38731 <= z3873_assgn38730;
        z3873_assgn38732 <= z3873_assgn38731;
        z3873_assgn38733 <= z3873_assgn38732;
        z3873_assgn38734 <= z3873_assgn38733;
        z3873_assgn38735 <= z3873_assgn38734;
        z3873_assgn38736 <= z3873_assgn38735;
        z3873_assgn38737 <= z3873_assgn38736;
        z3873_assgn38738 <= z3873_assgn38737;
        z3873_assgn38739 <= z3873_assgn38738;
        z3873_assgn387310 <= z3873_assgn38739;
        x8_G256_newbasis0 <= z3873_assgn387310;
        z4005_assgn40050 <= z4005_assgn4005;
        z4005_assgn40051 <= z4005_assgn40050;
        z4005_assgn40052 <= z4005_assgn40051;
        z4005_assgn40053 <= z4005_assgn40052;
        z4005_assgn40054 <= z4005_assgn40053;
        z4005_assgn40055 <= z4005_assgn40054;
        z4005_assgn40056 <= z4005_assgn40055;
        z4005_assgn40057 <= z4005_assgn40056;
        z4005_assgn40058 <= z4005_assgn40057;
        z4005_assgn40059 <= z4005_assgn40058;
        z4005_assgn400510 <= z4005_assgn40059;
        z_x8_G256_newbasis0 <= z4005_assgn400510;
        m0_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= m0_comar0_G4_mul0_G16_mul0_G256_inv0;
        m1_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= m1_comar0_G4_mul0_G16_mul0_G256_inv0;
        m3_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= m3_comar0_G4_mul0_G16_mul0_G256_inv0;
        m2_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= m2_comar0_G4_mul0_G16_mul0_G256_inv0;
        r0_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= r0_10_comar0_G4_mul0_G16_mul0_G256_inv0;
        r1_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= r1_10_comar0_G4_mul0_G16_mul0_G256_inv0;
        r2_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= r2_10_comar0_G4_mul0_G16_mul0_G256_inv0;
        r3_10_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= r3_10_comar0_G4_mul0_G16_mul0_G256_inv0;
        i1_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= i1_comar0_G4_mul0_G16_mul0_G256_inv0;
        i2_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= i2_comar0_G4_mul0_G16_mul0_G256_inv0;
        i0_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= i0_comar0_G4_mul0_G16_mul0_G256_inv0;
        i3_comar0_G4_mul0_G16_mul0_G256_inv0_reg <= i3_comar0_G4_mul0_G16_mul0_G256_inv0;
        e0_G4_mul0_G16_mul0_G256_inv0 <= (i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0);
        m0_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= m0_comar1_G4_mul0_G16_mul0_G256_inv0;
        m1_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= m1_comar1_G4_mul0_G16_mul0_G256_inv0;
        m3_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= m3_comar1_G4_mul0_G16_mul0_G256_inv0;
        m2_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= m2_comar1_G4_mul0_G16_mul0_G256_inv0;
        r0_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= r0_10_comar1_G4_mul0_G16_mul0_G256_inv0;
        r1_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= r1_10_comar1_G4_mul0_G16_mul0_G256_inv0;
        r2_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= r2_10_comar1_G4_mul0_G16_mul0_G256_inv0;
        r3_10_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= r3_10_comar1_G4_mul0_G16_mul0_G256_inv0;
        i1_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= i1_comar1_G4_mul0_G16_mul0_G256_inv0;
        i2_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= i2_comar1_G4_mul0_G16_mul0_G256_inv0;
        i0_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= i0_comar1_G4_mul0_G16_mul0_G256_inv0;
        i3_comar1_G4_mul0_G16_mul0_G256_inv0_reg <= i3_comar1_G4_mul0_G16_mul0_G256_inv0;
        p0_0_G4_mul0_G16_mul0_G256_inv0 <= (i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0);
        m0_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= m0_comar2_G4_mul0_G16_mul0_G256_inv0;
        m1_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= m1_comar2_G4_mul0_G16_mul0_G256_inv0;
        m3_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= m3_comar2_G4_mul0_G16_mul0_G256_inv0;
        m2_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= m2_comar2_G4_mul0_G16_mul0_G256_inv0;
        r0_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= r0_10_comar2_G4_mul0_G16_mul0_G256_inv0;
        r1_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= r1_10_comar2_G4_mul0_G16_mul0_G256_inv0;
        r2_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= r2_10_comar2_G4_mul0_G16_mul0_G256_inv0;
        r3_10_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= r3_10_comar2_G4_mul0_G16_mul0_G256_inv0;
        i1_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= i1_comar2_G4_mul0_G16_mul0_G256_inv0;
        i2_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= i2_comar2_G4_mul0_G16_mul0_G256_inv0;
        i0_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= i0_comar2_G4_mul0_G16_mul0_G256_inv0;
        i3_comar2_G4_mul0_G16_mul0_G256_inv0_reg <= i3_comar2_G4_mul0_G16_mul0_G256_inv0;
        q0_0_G4_mul0_G16_mul0_G256_inv0 <= (i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0);
        z4371_assgn43710 <= z4371_assgn4371;
        z4371_assgn43711 <= z4371_assgn43710;
        z691_assgn691 <= z4371_assgn43711;
        z4381_assgn43810 <= z4381_assgn4381;
        z4381_assgn43811 <= z4381_assgn43810;
        z699_assgn699 <= z4381_assgn43811;
        z4387_assgn43870 <= z4387_assgn4387;
        z4387_assgn43871 <= z4387_assgn43870;
        z703_assgn703 <= z4387_assgn43871;
        z4393_assgn43930 <= z4393_assgn4393;
        z4393_assgn43931 <= z4393_assgn43930;
        z707_assgn707 <= z4393_assgn43931;
        z4405_assgn44050 <= z4405_assgn4405;
        z4405_assgn44051 <= z4405_assgn44050;
        z717_assgn717 <= z4405_assgn44051;
        m0_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= m0_comar0_G4_mul1_G16_mul0_G256_inv0;
        m1_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= m1_comar0_G4_mul1_G16_mul0_G256_inv0;
        m3_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= m3_comar0_G4_mul1_G16_mul0_G256_inv0;
        m2_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= m2_comar0_G4_mul1_G16_mul0_G256_inv0;
        r0_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= r0_10_comar0_G4_mul1_G16_mul0_G256_inv0;
        r1_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= r1_10_comar0_G4_mul1_G16_mul0_G256_inv0;
        r2_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= r2_10_comar0_G4_mul1_G16_mul0_G256_inv0;
        r3_10_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= r3_10_comar0_G4_mul1_G16_mul0_G256_inv0;
        i1_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= i1_comar0_G4_mul1_G16_mul0_G256_inv0;
        i2_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= i2_comar0_G4_mul1_G16_mul0_G256_inv0;
        i0_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= i0_comar0_G4_mul1_G16_mul0_G256_inv0;
        i3_comar0_G4_mul1_G16_mul0_G256_inv0_reg <= i3_comar0_G4_mul1_G16_mul0_G256_inv0;
        e0_G4_mul1_G16_mul0_G256_inv0 <= (i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0);
        m0_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= m0_comar1_G4_mul1_G16_mul0_G256_inv0;
        m1_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= m1_comar1_G4_mul1_G16_mul0_G256_inv0;
        m3_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= m3_comar1_G4_mul1_G16_mul0_G256_inv0;
        m2_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= m2_comar1_G4_mul1_G16_mul0_G256_inv0;
        r0_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= r0_10_comar1_G4_mul1_G16_mul0_G256_inv0;
        r1_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= r1_10_comar1_G4_mul1_G16_mul0_G256_inv0;
        r2_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= r2_10_comar1_G4_mul1_G16_mul0_G256_inv0;
        r3_10_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= r3_10_comar1_G4_mul1_G16_mul0_G256_inv0;
        i1_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= i1_comar1_G4_mul1_G16_mul0_G256_inv0;
        i2_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= i2_comar1_G4_mul1_G16_mul0_G256_inv0;
        i0_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= i0_comar1_G4_mul1_G16_mul0_G256_inv0;
        i3_comar1_G4_mul1_G16_mul0_G256_inv0_reg <= i3_comar1_G4_mul1_G16_mul0_G256_inv0;
        p0_0_G4_mul1_G16_mul0_G256_inv0 <= (i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0);
        m0_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= m0_comar2_G4_mul1_G16_mul0_G256_inv0;
        m1_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= m1_comar2_G4_mul1_G16_mul0_G256_inv0;
        m3_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= m3_comar2_G4_mul1_G16_mul0_G256_inv0;
        m2_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= m2_comar2_G4_mul1_G16_mul0_G256_inv0;
        r0_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= r0_10_comar2_G4_mul1_G16_mul0_G256_inv0;
        r1_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= r1_10_comar2_G4_mul1_G16_mul0_G256_inv0;
        r2_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= r2_10_comar2_G4_mul1_G16_mul0_G256_inv0;
        r3_10_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= r3_10_comar2_G4_mul1_G16_mul0_G256_inv0;
        i1_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= i1_comar2_G4_mul1_G16_mul0_G256_inv0;
        i2_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= i2_comar2_G4_mul1_G16_mul0_G256_inv0;
        i0_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= i0_comar2_G4_mul1_G16_mul0_G256_inv0;
        i3_comar2_G4_mul1_G16_mul0_G256_inv0_reg <= i3_comar2_G4_mul1_G16_mul0_G256_inv0;
        q0_0_G4_mul1_G16_mul0_G256_inv0 <= (i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0);
        z4625_assgn46250 <= z4625_assgn4625;
        z4625_assgn46251 <= z4625_assgn46250;
        z935_assgn935 <= z4625_assgn46251;
        m0_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= m0_comar0_G4_mul2_G16_mul0_G256_inv0;
        m1_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= m1_comar0_G4_mul2_G16_mul0_G256_inv0;
        m3_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= m3_comar0_G4_mul2_G16_mul0_G256_inv0;
        m2_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= m2_comar0_G4_mul2_G16_mul0_G256_inv0;
        r0_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= r0_10_comar0_G4_mul2_G16_mul0_G256_inv0;
        r1_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= r1_10_comar0_G4_mul2_G16_mul0_G256_inv0;
        r2_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= r2_10_comar0_G4_mul2_G16_mul0_G256_inv0;
        r3_10_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= r3_10_comar0_G4_mul2_G16_mul0_G256_inv0;
        i1_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= i1_comar0_G4_mul2_G16_mul0_G256_inv0;
        i2_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= i2_comar0_G4_mul2_G16_mul0_G256_inv0;
        i0_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= i0_comar0_G4_mul2_G16_mul0_G256_inv0;
        i3_comar0_G4_mul2_G16_mul0_G256_inv0_reg <= i3_comar0_G4_mul2_G16_mul0_G256_inv0;
        e0_G4_mul2_G16_mul0_G256_inv0 <= (i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0);
        m0_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= m0_comar1_G4_mul2_G16_mul0_G256_inv0;
        m1_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= m1_comar1_G4_mul2_G16_mul0_G256_inv0;
        m3_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= m3_comar1_G4_mul2_G16_mul0_G256_inv0;
        m2_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= m2_comar1_G4_mul2_G16_mul0_G256_inv0;
        r0_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= r0_10_comar1_G4_mul2_G16_mul0_G256_inv0;
        r1_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= r1_10_comar1_G4_mul2_G16_mul0_G256_inv0;
        r2_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= r2_10_comar1_G4_mul2_G16_mul0_G256_inv0;
        r3_10_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= r3_10_comar1_G4_mul2_G16_mul0_G256_inv0;
        i1_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= i1_comar1_G4_mul2_G16_mul0_G256_inv0;
        i2_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= i2_comar1_G4_mul2_G16_mul0_G256_inv0;
        i0_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= i0_comar1_G4_mul2_G16_mul0_G256_inv0;
        i3_comar1_G4_mul2_G16_mul0_G256_inv0_reg <= i3_comar1_G4_mul2_G16_mul0_G256_inv0;
        p0_0_G4_mul2_G16_mul0_G256_inv0 <= (i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0);
        m0_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= m0_comar2_G4_mul2_G16_mul0_G256_inv0;
        m1_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= m1_comar2_G4_mul2_G16_mul0_G256_inv0;
        m3_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= m3_comar2_G4_mul2_G16_mul0_G256_inv0;
        m2_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= m2_comar2_G4_mul2_G16_mul0_G256_inv0;
        r0_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= r0_10_comar2_G4_mul2_G16_mul0_G256_inv0;
        r1_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= r1_10_comar2_G4_mul2_G16_mul0_G256_inv0;
        r2_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= r2_10_comar2_G4_mul2_G16_mul0_G256_inv0;
        r3_10_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= r3_10_comar2_G4_mul2_G16_mul0_G256_inv0;
        i1_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= i1_comar2_G4_mul2_G16_mul0_G256_inv0;
        i2_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= i2_comar2_G4_mul2_G16_mul0_G256_inv0;
        i0_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= i0_comar2_G4_mul2_G16_mul0_G256_inv0;
        i3_comar2_G4_mul2_G16_mul0_G256_inv0_reg <= i3_comar2_G4_mul2_G16_mul0_G256_inv0;
        q0_0_G4_mul2_G16_mul0_G256_inv0 <= (i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0);
        z4847_assgn48470 <= z4847_assgn4847;
        z4847_assgn48471 <= z4847_assgn48470;
        z1155_assgn1155 <= z4847_assgn48471;
        z4861_assgn48610 <= z4861_assgn4861;
        z4861_assgn48611 <= z4861_assgn48610;
        z1167_assgn1167 <= z4861_assgn48611;
        z4871_assgn48710 <= z4871_assgn4871;
        z4871_assgn48711 <= z4871_assgn48710;
        z1176_assgn1176 <= z4871_assgn48711;
        z4889_assgn48890 <= z4889_assgn4889;
        z4889_assgn48891 <= z4889_assgn48890;
        z1191_assgn1191 <= z4889_assgn48891;
        z4895_assgn48950 <= z4895_assgn4895;
        z4895_assgn48951 <= z4895_assgn48950;
        z1195_assgn1195 <= z4895_assgn48951;
        z4901_assgn49010 <= z4901_assgn4901;
        z4901_assgn49011 <= z4901_assgn49010;
        z1199_assgn1199 <= z4901_assgn49011;
        z4911_assgn49110 <= z4911_assgn4911;
        z4911_assgn49111 <= z4911_assgn49110;
        z1207_assgn1207 <= z4911_assgn49111;
        z4917_assgn49170 <= z4917_assgn4917;
        z4917_assgn49171 <= z4917_assgn49170;
        z1211_assgn1211 <= z4917_assgn49171;
        z4923_assgn49230 <= z4923_assgn4923;
        z4923_assgn49231 <= z4923_assgn49230;
        z1215_assgn1215 <= z4923_assgn49231;
        z4929_assgn49290 <= z4929_assgn4929;
        z4929_assgn49291 <= z4929_assgn49290;
        z1219_assgn1219 <= z4929_assgn49291;
        z4939_assgn49390 <= z4939_assgn4939;
        z4939_assgn49391 <= z4939_assgn49390;
        z1227_assgn1227 <= z4939_assgn49391;
        z4945_assgn49450 <= z4945_assgn4945;
        z4945_assgn49451 <= z4945_assgn49450;
        z1231_assgn1231 <= z4945_assgn49451;
        z4951_assgn49510 <= z4951_assgn4951;
        z4951_assgn49511 <= z4951_assgn49510;
        z1235_assgn1235 <= z4951_assgn49511;
        z4963_assgn49630 <= z4963_assgn4963;
        z4963_assgn49631 <= z4963_assgn49630;
        z1245_assgn1245 <= z4963_assgn49631;
        z4987_assgn49870 <= z4987_assgn4987;
        z4987_assgn49871 <= z4987_assgn49870;
        z1267_assgn1267 <= z4987_assgn49871;
        z4993_assgn49930 <= z4993_assgn4993;
        z4993_assgn49931 <= z4993_assgn49930;
        z1271_assgn1271 <= z4993_assgn49931;
        z4999_assgn49990 <= z4999_assgn4999;
        z4999_assgn49991 <= z4999_assgn49990;
        z1275_assgn1275 <= z4999_assgn49991;
        z5005_assgn50050 <= z5005_assgn5005;
        z5005_assgn50051 <= z5005_assgn50050;
        z1279_assgn1279 <= z5005_assgn50051;
        z5011_assgn50110 <= z5011_assgn5011;
        z5011_assgn50111 <= z5011_assgn50110;
        z1283_assgn1283 <= z5011_assgn50111;
        z5017_assgn50170 <= z5017_assgn5017;
        z5017_assgn50171 <= z5017_assgn50170;
        z1287_assgn1287 <= z5017_assgn50171;
        z5043_assgn50430 <= z5043_assgn5043;
        z5043_assgn50431 <= z5043_assgn50430;
        z1311_assgn1311 <= z5043_assgn50431;
        z5049_assgn50490 <= z5049_assgn5049;
        z5049_assgn50491 <= z5049_assgn50490;
        z1315_assgn1315 <= z5049_assgn50491;
        z5053_assgn50530 <= z5053_assgn5053;
        z5053_assgn50531 <= z5053_assgn50530;
        z5053_assgn50532 <= z5053_assgn50531;
        z1318_assgn1318 <= z5053_assgn50532;
        m1_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= m1_comar0_G4_mul3_G16_inv0_G256_inv0;
        z5057_assgn50570 <= z5057_assgn5057;
        z5057_assgn50571 <= z5057_assgn50570;
        z5057_assgn50572 <= z5057_assgn50571;
        z1319_assgn1319 <= z5057_assgn50572;
        m3_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= m3_comar0_G4_mul3_G16_inv0_G256_inv0;
        m0_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= m0_comar0_G4_mul3_G16_inv0_G256_inv0;
        m2_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= m2_comar0_G4_mul3_G16_inv0_G256_inv0;
        r0_10_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= r0_10_comar0_G4_mul3_G16_inv0_G256_inv0;
        z5067_assgn50670 <= z5067_assgn5067;
        z5067_assgn50671 <= z5067_assgn50670;
        z5067_assgn50672 <= z5067_assgn50671;
        z1327_assgn1327 <= z5067_assgn50672;
        z5071_assgn50710 <= z5071_assgn5071;
        z5071_assgn50711 <= z5071_assgn50710;
        z5071_assgn50712 <= z5071_assgn50711;
        z1329_assgn1329 <= z5071_assgn50712;
        z5075_assgn50750 <= z5075_assgn5075;
        z5075_assgn50751 <= z5075_assgn50750;
        z5075_assgn50752 <= z5075_assgn50751;
        z1331_assgn1331 <= z5075_assgn50752;
        i1_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= i1_comar0_G4_mul3_G16_inv0_G256_inv0;
        i2_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= i2_comar0_G4_mul3_G16_inv0_G256_inv0;
        z5081_assgn50810 <= z5081_assgn5081;
        z5081_assgn50811 <= z5081_assgn50810;
        z5081_assgn50812 <= z5081_assgn50811;
        z1336_assgn1336 <= z5081_assgn50812;
        i3_comar0_G4_mul3_G16_inv0_G256_inv0_reg <= i3_comar0_G4_mul3_G16_inv0_G256_inv0;
        e0_G4_mul3_G16_inv0_G256_inv0 <= (i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0);
        z5111_assgn51110 <= z5111_assgn5111;
        z5111_assgn51111 <= z5111_assgn51110;
        z1363_assgn1363 <= z5111_assgn51111;
        z5117_assgn51170 <= z5117_assgn5117;
        z5117_assgn51171 <= z5117_assgn51170;
        z1367_assgn1367 <= z5117_assgn51171;
        z5121_assgn51210 <= z5121_assgn5121;
        z5121_assgn51211 <= z5121_assgn51210;
        z5121_assgn51212 <= z5121_assgn51211;
        z1370_assgn1370 <= z5121_assgn51212;
        m1_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= m1_comar1_G4_mul3_G16_inv0_G256_inv0;
        z5125_assgn51250 <= z5125_assgn5125;
        z5125_assgn51251 <= z5125_assgn51250;
        z5125_assgn51252 <= z5125_assgn51251;
        z1371_assgn1371 <= z5125_assgn51252;
        m3_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= m3_comar1_G4_mul3_G16_inv0_G256_inv0;
        m0_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= m0_comar1_G4_mul3_G16_inv0_G256_inv0;
        m2_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= m2_comar1_G4_mul3_G16_inv0_G256_inv0;
        r0_10_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= r0_10_comar1_G4_mul3_G16_inv0_G256_inv0;
        z5135_assgn51350 <= z5135_assgn5135;
        z5135_assgn51351 <= z5135_assgn51350;
        z5135_assgn51352 <= z5135_assgn51351;
        z1379_assgn1379 <= z5135_assgn51352;
        z5139_assgn51390 <= z5139_assgn5139;
        z5139_assgn51391 <= z5139_assgn51390;
        z5139_assgn51392 <= z5139_assgn51391;
        z1381_assgn1381 <= z5139_assgn51392;
        z5143_assgn51430 <= z5143_assgn5143;
        z5143_assgn51431 <= z5143_assgn51430;
        z5143_assgn51432 <= z5143_assgn51431;
        z1383_assgn1383 <= z5143_assgn51432;
        i1_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= i1_comar1_G4_mul3_G16_inv0_G256_inv0;
        i2_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= i2_comar1_G4_mul3_G16_inv0_G256_inv0;
        z5149_assgn51490 <= z5149_assgn5149;
        z5149_assgn51491 <= z5149_assgn51490;
        z5149_assgn51492 <= z5149_assgn51491;
        z1388_assgn1388 <= z5149_assgn51492;
        i3_comar1_G4_mul3_G16_inv0_G256_inv0_reg <= i3_comar1_G4_mul3_G16_inv0_G256_inv0;
        p0_0_G4_mul3_G16_inv0_G256_inv0 <= (i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0);
        z5183_assgn51830 <= z5183_assgn5183;
        z5183_assgn51831 <= z5183_assgn51830;
        z1419_assgn1419 <= z5183_assgn51831;
        z5189_assgn51890 <= z5189_assgn5189;
        z5189_assgn51891 <= z5189_assgn51890;
        z1423_assgn1423 <= z5189_assgn51891;
        z5193_assgn51930 <= z5193_assgn5193;
        z5193_assgn51931 <= z5193_assgn51930;
        z5193_assgn51932 <= z5193_assgn51931;
        z1426_assgn1426 <= z5193_assgn51932;
        m1_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= m1_comar2_G4_mul3_G16_inv0_G256_inv0;
        z5197_assgn51970 <= z5197_assgn5197;
        z5197_assgn51971 <= z5197_assgn51970;
        z5197_assgn51972 <= z5197_assgn51971;
        z1427_assgn1427 <= z5197_assgn51972;
        m3_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= m3_comar2_G4_mul3_G16_inv0_G256_inv0;
        m0_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= m0_comar2_G4_mul3_G16_inv0_G256_inv0;
        m2_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= m2_comar2_G4_mul3_G16_inv0_G256_inv0;
        r0_10_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= r0_10_comar2_G4_mul3_G16_inv0_G256_inv0;
        z5207_assgn52070 <= z5207_assgn5207;
        z5207_assgn52071 <= z5207_assgn52070;
        z5207_assgn52072 <= z5207_assgn52071;
        z1435_assgn1435 <= z5207_assgn52072;
        z5211_assgn52110 <= z5211_assgn5211;
        z5211_assgn52111 <= z5211_assgn52110;
        z5211_assgn52112 <= z5211_assgn52111;
        z1437_assgn1437 <= z5211_assgn52112;
        z5215_assgn52150 <= z5215_assgn5215;
        z5215_assgn52151 <= z5215_assgn52150;
        z5215_assgn52152 <= z5215_assgn52151;
        z1439_assgn1439 <= z5215_assgn52152;
        i1_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= i1_comar2_G4_mul3_G16_inv0_G256_inv0;
        i2_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= i2_comar2_G4_mul3_G16_inv0_G256_inv0;
        z5221_assgn52210 <= z5221_assgn5221;
        z5221_assgn52211 <= z5221_assgn52210;
        z5221_assgn52212 <= z5221_assgn52211;
        z1444_assgn1444 <= z5221_assgn52212;
        i3_comar2_G4_mul3_G16_inv0_G256_inv0_reg <= i3_comar2_G4_mul3_G16_inv0_G256_inv0;
        q0_0_G4_mul3_G16_inv0_G256_inv0 <= (i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0);
        z5243_assgn52430 <= z5243_assgn5243;
        z5243_assgn52431 <= z5243_assgn52430;
        z5243_assgn52432 <= z5243_assgn52431;
        z5243_assgn52433 <= z5243_assgn52432;
        z5243_assgn52434 <= z5243_assgn52433;
        z1463_assgn1463 <= z5243_assgn52434;
        z5253_assgn52530 <= z5253_assgn5253;
        z5253_assgn52531 <= z5253_assgn52530;
        z1472_assgn1472 <= z5253_assgn52531;
        z5259_assgn52590 <= z5259_assgn5259;
        z5259_assgn52591 <= z5259_assgn52590;
        z5259_assgn52592 <= z5259_assgn52591;
        z5259_assgn52593 <= z5259_assgn52592;
        z5259_assgn52594 <= z5259_assgn52593;
        z1475_assgn1475 <= z5259_assgn52594;
        z5265_assgn52650 <= z5265_assgn5265;
        z5265_assgn52651 <= z5265_assgn52650;
        z5265_assgn52652 <= z5265_assgn52651;
        z5265_assgn52653 <= z5265_assgn52652;
        z5265_assgn52654 <= z5265_assgn52653;
        z1479_assgn1479 <= z5265_assgn52654;
        z5271_assgn52710 <= z5271_assgn5271;
        z5271_assgn52711 <= z5271_assgn52710;
        z5271_assgn52712 <= z5271_assgn52711;
        z5271_assgn52713 <= z5271_assgn52712;
        z5271_assgn52714 <= z5271_assgn52713;
        z1483_assgn1483 <= z5271_assgn52714;
        z5277_assgn52770 <= z5277_assgn5277;
        z5277_assgn52771 <= z5277_assgn52770;
        z5277_assgn52772 <= z5277_assgn52771;
        z5277_assgn52773 <= z5277_assgn52772;
        z5277_assgn52774 <= z5277_assgn52773;
        z1487_assgn1487 <= z5277_assgn52774;
        z5299_assgn52990 <= z5299_assgn5299;
        z5299_assgn52991 <= z5299_assgn52990;
        z5299_assgn52992 <= z5299_assgn52991;
        z5299_assgn52993 <= z5299_assgn52992;
        z5299_assgn52994 <= z5299_assgn52993;
        z1507_assgn1507 <= z5299_assgn52994;
        z5305_assgn53050 <= z5305_assgn5305;
        z5305_assgn53051 <= z5305_assgn53050;
        z5305_assgn53052 <= z5305_assgn53051;
        z5305_assgn53053 <= z5305_assgn53052;
        z5305_assgn53054 <= z5305_assgn53053;
        z1511_assgn1511 <= z5305_assgn53054;
        z5311_assgn53110 <= z5311_assgn5311;
        z5311_assgn53111 <= z5311_assgn53110;
        z5311_assgn53112 <= z5311_assgn53111;
        z5311_assgn53113 <= z5311_assgn53112;
        z5311_assgn53114 <= z5311_assgn53113;
        z1515_assgn1515 <= z5311_assgn53114;
        z5317_assgn53170 <= z5317_assgn5317;
        z5317_assgn53171 <= z5317_assgn53170;
        z1519_assgn1519 <= z5317_assgn53171;
        z5323_assgn53230 <= z5323_assgn5323;
        z5323_assgn53231 <= z5323_assgn53230;
        z1523_assgn1523 <= z5323_assgn53231;
        z5329_assgn53290 <= z5329_assgn5329;
        z5329_assgn53291 <= z5329_assgn53290;
        z1527_assgn1527 <= z5329_assgn53291;
        z5355_assgn53550 <= z5355_assgn5355;
        z5355_assgn53551 <= z5355_assgn53550;
        z1551_assgn1551 <= z5355_assgn53551;
        z5361_assgn53610 <= z5361_assgn5361;
        z5361_assgn53611 <= z5361_assgn53610;
        z5361_assgn53612 <= z5361_assgn53611;
        z5361_assgn53613 <= z5361_assgn53612;
        z5361_assgn53614 <= z5361_assgn53613;
        z1555_assgn1555 <= z5361_assgn53614;
        z5365_assgn53650 <= z5365_assgn5365;
        z5365_assgn53651 <= z5365_assgn53650;
        z5365_assgn53652 <= z5365_assgn53651;
        z1558_assgn1558 <= z5365_assgn53652;
        m1_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= m1_comar0_G4_mul4_G16_inv0_G256_inv0;
        z5369_assgn53690 <= z5369_assgn5369;
        z5369_assgn53691 <= z5369_assgn53690;
        z5369_assgn53692 <= z5369_assgn53691;
        z5369_assgn53693 <= z5369_assgn53692;
        z5369_assgn53694 <= z5369_assgn53693;
        z5369_assgn53695 <= z5369_assgn53694;
        z1559_assgn1559 <= z5369_assgn53695;
        m3_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= m3_comar0_G4_mul4_G16_inv0_G256_inv0;
        m0_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= m0_comar0_G4_mul4_G16_inv0_G256_inv0;
        m2_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= m2_comar0_G4_mul4_G16_inv0_G256_inv0;
        z5375_assgn53750 <= z5375_assgn5375;
        z5375_assgn53751 <= z5375_assgn53750;
        z5375_assgn53752 <= z5375_assgn53751;
        z1563_assgn1563 <= z5375_assgn53752;
        r0_10_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= r0_10_comar0_G4_mul4_G16_inv0_G256_inv0;
        z5381_assgn53810 <= z5381_assgn5381;
        z5381_assgn53811 <= z5381_assgn53810;
        z5381_assgn53812 <= z5381_assgn53811;
        z1567_assgn1567 <= z5381_assgn53812;
        z5385_assgn53850 <= z5385_assgn5385;
        z5385_assgn53851 <= z5385_assgn53850;
        z5385_assgn53852 <= z5385_assgn53851;
        z5385_assgn53853 <= z5385_assgn53852;
        z5385_assgn53854 <= z5385_assgn53853;
        z5385_assgn53855 <= z5385_assgn53854;
        z1569_assgn1569 <= z5385_assgn53855;
        z5389_assgn53890 <= z5389_assgn5389;
        z5389_assgn53891 <= z5389_assgn53890;
        z5389_assgn53892 <= z5389_assgn53891;
        z5389_assgn53893 <= z5389_assgn53892;
        z5389_assgn53894 <= z5389_assgn53893;
        z5389_assgn53895 <= z5389_assgn53894;
        z1571_assgn1571 <= z5389_assgn53895;
        z5393_assgn53930 <= z5393_assgn5393;
        z5393_assgn53931 <= z5393_assgn53930;
        z5393_assgn53932 <= z5393_assgn53931;
        z1574_assgn1574 <= z5393_assgn53932;
        i2_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= i2_comar0_G4_mul4_G16_inv0_G256_inv0;
        z5397_assgn53970 <= z5397_assgn5397;
        z5397_assgn53971 <= z5397_assgn53970;
        z5397_assgn53972 <= z5397_assgn53971;
        z5397_assgn53973 <= z5397_assgn53972;
        z5397_assgn53974 <= z5397_assgn53973;
        z5397_assgn53975 <= z5397_assgn53974;
        z1576_assgn1576 <= z5397_assgn53975;
        i3_comar0_G4_mul4_G16_inv0_G256_inv0_reg <= i3_comar0_G4_mul4_G16_inv0_G256_inv0;
        e0_G4_mul4_G16_inv0_G256_inv0 <= (i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0);
        z5427_assgn54270 <= z5427_assgn5427;
        z5427_assgn54271 <= z5427_assgn54270;
        z1603_assgn1603 <= z5427_assgn54271;
        z5433_assgn54330 <= z5433_assgn5433;
        z5433_assgn54331 <= z5433_assgn54330;
        z5433_assgn54332 <= z5433_assgn54331;
        z5433_assgn54333 <= z5433_assgn54332;
        z5433_assgn54334 <= z5433_assgn54333;
        z1607_assgn1607 <= z5433_assgn54334;
        z5437_assgn54370 <= z5437_assgn5437;
        z5437_assgn54371 <= z5437_assgn54370;
        z5437_assgn54372 <= z5437_assgn54371;
        z1610_assgn1610 <= z5437_assgn54372;
        m1_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= m1_comar1_G4_mul4_G16_inv0_G256_inv0;
        z5441_assgn54410 <= z5441_assgn5441;
        z5441_assgn54411 <= z5441_assgn54410;
        z5441_assgn54412 <= z5441_assgn54411;
        z5441_assgn54413 <= z5441_assgn54412;
        z5441_assgn54414 <= z5441_assgn54413;
        z5441_assgn54415 <= z5441_assgn54414;
        z1611_assgn1611 <= z5441_assgn54415;
        m3_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= m3_comar1_G4_mul4_G16_inv0_G256_inv0;
        m0_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= m0_comar1_G4_mul4_G16_inv0_G256_inv0;
        m2_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= m2_comar1_G4_mul4_G16_inv0_G256_inv0;
        z5447_assgn54470 <= z5447_assgn5447;
        z5447_assgn54471 <= z5447_assgn54470;
        z5447_assgn54472 <= z5447_assgn54471;
        z1615_assgn1615 <= z5447_assgn54472;
        r0_10_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= r0_10_comar1_G4_mul4_G16_inv0_G256_inv0;
        z5453_assgn54530 <= z5453_assgn5453;
        z5453_assgn54531 <= z5453_assgn54530;
        z5453_assgn54532 <= z5453_assgn54531;
        z1619_assgn1619 <= z5453_assgn54532;
        z5457_assgn54570 <= z5457_assgn5457;
        z5457_assgn54571 <= z5457_assgn54570;
        z5457_assgn54572 <= z5457_assgn54571;
        z5457_assgn54573 <= z5457_assgn54572;
        z5457_assgn54574 <= z5457_assgn54573;
        z5457_assgn54575 <= z5457_assgn54574;
        z1621_assgn1621 <= z5457_assgn54575;
        z5461_assgn54610 <= z5461_assgn5461;
        z5461_assgn54611 <= z5461_assgn54610;
        z5461_assgn54612 <= z5461_assgn54611;
        z5461_assgn54613 <= z5461_assgn54612;
        z5461_assgn54614 <= z5461_assgn54613;
        z5461_assgn54615 <= z5461_assgn54614;
        z1623_assgn1623 <= z5461_assgn54615;
        z5465_assgn54650 <= z5465_assgn5465;
        z5465_assgn54651 <= z5465_assgn54650;
        z5465_assgn54652 <= z5465_assgn54651;
        z1626_assgn1626 <= z5465_assgn54652;
        i2_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= i2_comar1_G4_mul4_G16_inv0_G256_inv0;
        z5469_assgn54690 <= z5469_assgn5469;
        z5469_assgn54691 <= z5469_assgn54690;
        z5469_assgn54692 <= z5469_assgn54691;
        z5469_assgn54693 <= z5469_assgn54692;
        z5469_assgn54694 <= z5469_assgn54693;
        z5469_assgn54695 <= z5469_assgn54694;
        z1628_assgn1628 <= z5469_assgn54695;
        i3_comar1_G4_mul4_G16_inv0_G256_inv0_reg <= i3_comar1_G4_mul4_G16_inv0_G256_inv0;
        p0_0_G4_mul4_G16_inv0_G256_inv0 <= (i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0);
        z5503_assgn55030 <= z5503_assgn5503;
        z5503_assgn55031 <= z5503_assgn55030;
        z1659_assgn1659 <= z5503_assgn55031;
        z5509_assgn55090 <= z5509_assgn5509;
        z5509_assgn55091 <= z5509_assgn55090;
        z5509_assgn55092 <= z5509_assgn55091;
        z5509_assgn55093 <= z5509_assgn55092;
        z5509_assgn55094 <= z5509_assgn55093;
        z1663_assgn1663 <= z5509_assgn55094;
        z5513_assgn55130 <= z5513_assgn5513;
        z5513_assgn55131 <= z5513_assgn55130;
        z5513_assgn55132 <= z5513_assgn55131;
        z1666_assgn1666 <= z5513_assgn55132;
        m1_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= m1_comar2_G4_mul4_G16_inv0_G256_inv0;
        z5517_assgn55170 <= z5517_assgn5517;
        z5517_assgn55171 <= z5517_assgn55170;
        z5517_assgn55172 <= z5517_assgn55171;
        z5517_assgn55173 <= z5517_assgn55172;
        z5517_assgn55174 <= z5517_assgn55173;
        z5517_assgn55175 <= z5517_assgn55174;
        z1667_assgn1667 <= z5517_assgn55175;
        m3_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= m3_comar2_G4_mul4_G16_inv0_G256_inv0;
        m0_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= m0_comar2_G4_mul4_G16_inv0_G256_inv0;
        m2_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= m2_comar2_G4_mul4_G16_inv0_G256_inv0;
        z5523_assgn55230 <= z5523_assgn5523;
        z5523_assgn55231 <= z5523_assgn55230;
        z5523_assgn55232 <= z5523_assgn55231;
        z1671_assgn1671 <= z5523_assgn55232;
        r0_10_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= r0_10_comar2_G4_mul4_G16_inv0_G256_inv0;
        z5529_assgn55290 <= z5529_assgn5529;
        z5529_assgn55291 <= z5529_assgn55290;
        z5529_assgn55292 <= z5529_assgn55291;
        z1675_assgn1675 <= z5529_assgn55292;
        z5533_assgn55330 <= z5533_assgn5533;
        z5533_assgn55331 <= z5533_assgn55330;
        z5533_assgn55332 <= z5533_assgn55331;
        z5533_assgn55333 <= z5533_assgn55332;
        z5533_assgn55334 <= z5533_assgn55333;
        z5533_assgn55335 <= z5533_assgn55334;
        z1677_assgn1677 <= z5533_assgn55335;
        z5537_assgn55370 <= z5537_assgn5537;
        z5537_assgn55371 <= z5537_assgn55370;
        z5537_assgn55372 <= z5537_assgn55371;
        z5537_assgn55373 <= z5537_assgn55372;
        z5537_assgn55374 <= z5537_assgn55373;
        z5537_assgn55375 <= z5537_assgn55374;
        z1679_assgn1679 <= z5537_assgn55375;
        z5541_assgn55410 <= z5541_assgn5541;
        z5541_assgn55411 <= z5541_assgn55410;
        z5541_assgn55412 <= z5541_assgn55411;
        z1682_assgn1682 <= z5541_assgn55412;
        i2_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= i2_comar2_G4_mul4_G16_inv0_G256_inv0;
        z5545_assgn55450 <= z5545_assgn5545;
        z5545_assgn55451 <= z5545_assgn55450;
        z5545_assgn55452 <= z5545_assgn55451;
        z5545_assgn55453 <= z5545_assgn55452;
        z5545_assgn55454 <= z5545_assgn55453;
        z5545_assgn55455 <= z5545_assgn55454;
        z1684_assgn1684 <= z5545_assgn55455;
        i3_comar2_G4_mul4_G16_inv0_G256_inv0_reg <= i3_comar2_G4_mul4_G16_inv0_G256_inv0;
        q0_0_G4_mul4_G16_inv0_G256_inv0 <= (i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0);
        z5567_assgn55670 <= z5567_assgn5567;
        z5567_assgn55671 <= z5567_assgn55670;
        z5567_assgn55672 <= z5567_assgn55671;
        z5567_assgn55673 <= z5567_assgn55672;
        z5567_assgn55674 <= z5567_assgn55673;
        z5567_assgn55675 <= z5567_assgn55674;
        z5567_assgn55676 <= z5567_assgn55675;
        z5567_assgn55677 <= z5567_assgn55676;
        z1703_assgn1703 <= z5567_assgn55677;
        z5589_assgn55890 <= z5589_assgn5589;
        z5589_assgn55891 <= z5589_assgn55890;
        z5589_assgn55892 <= z5589_assgn55891;
        z5589_assgn55893 <= z5589_assgn55892;
        z5589_assgn55894 <= z5589_assgn55893;
        z1723_assgn1723 <= z5589_assgn55894;
        z5595_assgn55950 <= z5595_assgn5595;
        z5595_assgn55951 <= z5595_assgn55950;
        z5595_assgn55952 <= z5595_assgn55951;
        z5595_assgn55953 <= z5595_assgn55952;
        z5595_assgn55954 <= z5595_assgn55953;
        z1727_assgn1727 <= z5595_assgn55954;
        z5601_assgn56010 <= z5601_assgn5601;
        z5601_assgn56011 <= z5601_assgn56010;
        z5601_assgn56012 <= z5601_assgn56011;
        z5601_assgn56013 <= z5601_assgn56012;
        z5601_assgn56014 <= z5601_assgn56013;
        z1731_assgn1731 <= z5601_assgn56014;
        z5607_assgn56070 <= z5607_assgn5607;
        z5607_assgn56071 <= z5607_assgn56070;
        z1735_assgn1735 <= z5607_assgn56071;
        z5613_assgn56130 <= z5613_assgn5613;
        z5613_assgn56131 <= z5613_assgn56130;
        z1739_assgn1739 <= z5613_assgn56131;
        z5619_assgn56190 <= z5619_assgn5619;
        z5619_assgn56191 <= z5619_assgn56190;
        z1743_assgn1743 <= z5619_assgn56191;
        z5645_assgn56450 <= z5645_assgn5645;
        z5645_assgn56451 <= z5645_assgn56450;
        z1767_assgn1767 <= z5645_assgn56451;
        z5651_assgn56510 <= z5651_assgn5651;
        z5651_assgn56511 <= z5651_assgn56510;
        z5651_assgn56512 <= z5651_assgn56511;
        z5651_assgn56513 <= z5651_assgn56512;
        z5651_assgn56514 <= z5651_assgn56513;
        z1771_assgn1771 <= z5651_assgn56514;
        z5655_assgn56550 <= z5655_assgn5655;
        z5655_assgn56551 <= z5655_assgn56550;
        z5655_assgn56552 <= z5655_assgn56551;
        z1774_assgn1774 <= z5655_assgn56552;
        m1_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= m1_comar0_G4_mul5_G16_inv0_G256_inv0;
        z5659_assgn56590 <= z5659_assgn5659;
        z5659_assgn56591 <= z5659_assgn56590;
        z5659_assgn56592 <= z5659_assgn56591;
        z5659_assgn56593 <= z5659_assgn56592;
        z5659_assgn56594 <= z5659_assgn56593;
        z5659_assgn56595 <= z5659_assgn56594;
        z1775_assgn1775 <= z5659_assgn56595;
        m3_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= m3_comar0_G4_mul5_G16_inv0_G256_inv0;
        m0_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= m0_comar0_G4_mul5_G16_inv0_G256_inv0;
        m2_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= m2_comar0_G4_mul5_G16_inv0_G256_inv0;
        z5665_assgn56650 <= z5665_assgn5665;
        z5665_assgn56651 <= z5665_assgn56650;
        z5665_assgn56652 <= z5665_assgn56651;
        z1779_assgn1779 <= z5665_assgn56652;
        r0_10_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= r0_10_comar0_G4_mul5_G16_inv0_G256_inv0;
        z5671_assgn56710 <= z5671_assgn5671;
        z5671_assgn56711 <= z5671_assgn56710;
        z5671_assgn56712 <= z5671_assgn56711;
        z1783_assgn1783 <= z5671_assgn56712;
        z5675_assgn56750 <= z5675_assgn5675;
        z5675_assgn56751 <= z5675_assgn56750;
        z5675_assgn56752 <= z5675_assgn56751;
        z5675_assgn56753 <= z5675_assgn56752;
        z5675_assgn56754 <= z5675_assgn56753;
        z5675_assgn56755 <= z5675_assgn56754;
        z1785_assgn1785 <= z5675_assgn56755;
        z5679_assgn56790 <= z5679_assgn5679;
        z5679_assgn56791 <= z5679_assgn56790;
        z5679_assgn56792 <= z5679_assgn56791;
        z5679_assgn56793 <= z5679_assgn56792;
        z5679_assgn56794 <= z5679_assgn56793;
        z5679_assgn56795 <= z5679_assgn56794;
        z1787_assgn1787 <= z5679_assgn56795;
        z5683_assgn56830 <= z5683_assgn5683;
        z5683_assgn56831 <= z5683_assgn56830;
        z5683_assgn56832 <= z5683_assgn56831;
        z1790_assgn1790 <= z5683_assgn56832;
        i2_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= i2_comar0_G4_mul5_G16_inv0_G256_inv0;
        z5687_assgn56870 <= z5687_assgn5687;
        z5687_assgn56871 <= z5687_assgn56870;
        z5687_assgn56872 <= z5687_assgn56871;
        z5687_assgn56873 <= z5687_assgn56872;
        z5687_assgn56874 <= z5687_assgn56873;
        z5687_assgn56875 <= z5687_assgn56874;
        z1792_assgn1792 <= z5687_assgn56875;
        i3_comar0_G4_mul5_G16_inv0_G256_inv0_reg <= i3_comar0_G4_mul5_G16_inv0_G256_inv0;
        e0_G4_mul5_G16_inv0_G256_inv0 <= (i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0);
        z5717_assgn57170 <= z5717_assgn5717;
        z5717_assgn57171 <= z5717_assgn57170;
        z1819_assgn1819 <= z5717_assgn57171;
        z5723_assgn57230 <= z5723_assgn5723;
        z5723_assgn57231 <= z5723_assgn57230;
        z5723_assgn57232 <= z5723_assgn57231;
        z5723_assgn57233 <= z5723_assgn57232;
        z5723_assgn57234 <= z5723_assgn57233;
        z1823_assgn1823 <= z5723_assgn57234;
        z5727_assgn57270 <= z5727_assgn5727;
        z5727_assgn57271 <= z5727_assgn57270;
        z5727_assgn57272 <= z5727_assgn57271;
        z1826_assgn1826 <= z5727_assgn57272;
        m1_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= m1_comar1_G4_mul5_G16_inv0_G256_inv0;
        z5731_assgn57310 <= z5731_assgn5731;
        z5731_assgn57311 <= z5731_assgn57310;
        z5731_assgn57312 <= z5731_assgn57311;
        z5731_assgn57313 <= z5731_assgn57312;
        z5731_assgn57314 <= z5731_assgn57313;
        z5731_assgn57315 <= z5731_assgn57314;
        z1827_assgn1827 <= z5731_assgn57315;
        m3_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= m3_comar1_G4_mul5_G16_inv0_G256_inv0;
        m0_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= m0_comar1_G4_mul5_G16_inv0_G256_inv0;
        m2_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= m2_comar1_G4_mul5_G16_inv0_G256_inv0;
        z5737_assgn57370 <= z5737_assgn5737;
        z5737_assgn57371 <= z5737_assgn57370;
        z5737_assgn57372 <= z5737_assgn57371;
        z1831_assgn1831 <= z5737_assgn57372;
        r0_10_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= r0_10_comar1_G4_mul5_G16_inv0_G256_inv0;
        z5743_assgn57430 <= z5743_assgn5743;
        z5743_assgn57431 <= z5743_assgn57430;
        z5743_assgn57432 <= z5743_assgn57431;
        z1835_assgn1835 <= z5743_assgn57432;
        z5747_assgn57470 <= z5747_assgn5747;
        z5747_assgn57471 <= z5747_assgn57470;
        z5747_assgn57472 <= z5747_assgn57471;
        z5747_assgn57473 <= z5747_assgn57472;
        z5747_assgn57474 <= z5747_assgn57473;
        z5747_assgn57475 <= z5747_assgn57474;
        z1837_assgn1837 <= z5747_assgn57475;
        z5751_assgn57510 <= z5751_assgn5751;
        z5751_assgn57511 <= z5751_assgn57510;
        z5751_assgn57512 <= z5751_assgn57511;
        z5751_assgn57513 <= z5751_assgn57512;
        z5751_assgn57514 <= z5751_assgn57513;
        z5751_assgn57515 <= z5751_assgn57514;
        z1839_assgn1839 <= z5751_assgn57515;
        z5755_assgn57550 <= z5755_assgn5755;
        z5755_assgn57551 <= z5755_assgn57550;
        z5755_assgn57552 <= z5755_assgn57551;
        z1842_assgn1842 <= z5755_assgn57552;
        i2_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= i2_comar1_G4_mul5_G16_inv0_G256_inv0;
        z5759_assgn57590 <= z5759_assgn5759;
        z5759_assgn57591 <= z5759_assgn57590;
        z5759_assgn57592 <= z5759_assgn57591;
        z5759_assgn57593 <= z5759_assgn57592;
        z5759_assgn57594 <= z5759_assgn57593;
        z5759_assgn57595 <= z5759_assgn57594;
        z1844_assgn1844 <= z5759_assgn57595;
        i3_comar1_G4_mul5_G16_inv0_G256_inv0_reg <= i3_comar1_G4_mul5_G16_inv0_G256_inv0;
        p0_0_G4_mul5_G16_inv0_G256_inv0 <= (i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0);
        z5793_assgn57930 <= z5793_assgn5793;
        z5793_assgn57931 <= z5793_assgn57930;
        z1875_assgn1875 <= z5793_assgn57931;
        z5799_assgn57990 <= z5799_assgn5799;
        z5799_assgn57991 <= z5799_assgn57990;
        z5799_assgn57992 <= z5799_assgn57991;
        z5799_assgn57993 <= z5799_assgn57992;
        z5799_assgn57994 <= z5799_assgn57993;
        z1879_assgn1879 <= z5799_assgn57994;
        z5803_assgn58030 <= z5803_assgn5803;
        z5803_assgn58031 <= z5803_assgn58030;
        z5803_assgn58032 <= z5803_assgn58031;
        z1882_assgn1882 <= z5803_assgn58032;
        m1_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= m1_comar2_G4_mul5_G16_inv0_G256_inv0;
        z5807_assgn58070 <= z5807_assgn5807;
        z5807_assgn58071 <= z5807_assgn58070;
        z5807_assgn58072 <= z5807_assgn58071;
        z5807_assgn58073 <= z5807_assgn58072;
        z5807_assgn58074 <= z5807_assgn58073;
        z5807_assgn58075 <= z5807_assgn58074;
        z1883_assgn1883 <= z5807_assgn58075;
        m3_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= m3_comar2_G4_mul5_G16_inv0_G256_inv0;
        m0_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= m0_comar2_G4_mul5_G16_inv0_G256_inv0;
        m2_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= m2_comar2_G4_mul5_G16_inv0_G256_inv0;
        z5813_assgn58130 <= z5813_assgn5813;
        z5813_assgn58131 <= z5813_assgn58130;
        z5813_assgn58132 <= z5813_assgn58131;
        z1887_assgn1887 <= z5813_assgn58132;
        r0_10_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= r0_10_comar2_G4_mul5_G16_inv0_G256_inv0;
        z5819_assgn58190 <= z5819_assgn5819;
        z5819_assgn58191 <= z5819_assgn58190;
        z5819_assgn58192 <= z5819_assgn58191;
        z1891_assgn1891 <= z5819_assgn58192;
        z5823_assgn58230 <= z5823_assgn5823;
        z5823_assgn58231 <= z5823_assgn58230;
        z5823_assgn58232 <= z5823_assgn58231;
        z5823_assgn58233 <= z5823_assgn58232;
        z5823_assgn58234 <= z5823_assgn58233;
        z5823_assgn58235 <= z5823_assgn58234;
        z1893_assgn1893 <= z5823_assgn58235;
        z5827_assgn58270 <= z5827_assgn5827;
        z5827_assgn58271 <= z5827_assgn58270;
        z5827_assgn58272 <= z5827_assgn58271;
        z5827_assgn58273 <= z5827_assgn58272;
        z5827_assgn58274 <= z5827_assgn58273;
        z5827_assgn58275 <= z5827_assgn58274;
        z1895_assgn1895 <= z5827_assgn58275;
        z5831_assgn58310 <= z5831_assgn5831;
        z5831_assgn58311 <= z5831_assgn58310;
        z5831_assgn58312 <= z5831_assgn58311;
        z1898_assgn1898 <= z5831_assgn58312;
        i2_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= i2_comar2_G4_mul5_G16_inv0_G256_inv0;
        z5835_assgn58350 <= z5835_assgn5835;
        z5835_assgn58351 <= z5835_assgn58350;
        z5835_assgn58352 <= z5835_assgn58351;
        z5835_assgn58353 <= z5835_assgn58352;
        z5835_assgn58354 <= z5835_assgn58353;
        z5835_assgn58355 <= z5835_assgn58354;
        z1900_assgn1900 <= z5835_assgn58355;
        i3_comar2_G4_mul5_G16_inv0_G256_inv0_reg <= i3_comar2_G4_mul5_G16_inv0_G256_inv0;
        q0_0_G4_mul5_G16_inv0_G256_inv0 <= (i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0);
        z5857_assgn58570 <= z5857_assgn5857;
        z5857_assgn58571 <= z5857_assgn58570;
        z5857_assgn58572 <= z5857_assgn58571;
        z5857_assgn58573 <= z5857_assgn58572;
        z5857_assgn58574 <= z5857_assgn58573;
        z5857_assgn58575 <= z5857_assgn58574;
        z5857_assgn58576 <= z5857_assgn58575;
        z5857_assgn58577 <= z5857_assgn58576;
        z1919_assgn1919 <= z5857_assgn58577;
        z5867_assgn58670 <= z5867_assgn5867;
        z5867_assgn58671 <= z5867_assgn58670;
        z5867_assgn58672 <= z5867_assgn58671;
        z5867_assgn58673 <= z5867_assgn58672;
        z5867_assgn58674 <= z5867_assgn58673;
        z5867_assgn58675 <= z5867_assgn58674;
        z5867_assgn58676 <= z5867_assgn58675;
        z5867_assgn58677 <= z5867_assgn58676;
        z1927_assgn1927 <= z5867_assgn58677;
        z5889_assgn58890 <= z5889_assgn5889;
        z5889_assgn58891 <= z5889_assgn58890;
        z5889_assgn58892 <= z5889_assgn58891;
        z5889_assgn58893 <= z5889_assgn58892;
        z5889_assgn58894 <= z5889_assgn58893;
        z5889_assgn58895 <= z5889_assgn58894;
        z5889_assgn58896 <= z5889_assgn58895;
        z5889_assgn58897 <= z5889_assgn58896;
        z1947_assgn1947 <= z5889_assgn58897;
        z5895_assgn58950 <= z5895_assgn5895;
        z5895_assgn58951 <= z5895_assgn58950;
        z5895_assgn58952 <= z5895_assgn58951;
        z5895_assgn58953 <= z5895_assgn58952;
        z5895_assgn58954 <= z5895_assgn58953;
        z5895_assgn58955 <= z5895_assgn58954;
        z5895_assgn58956 <= z5895_assgn58955;
        z5895_assgn58957 <= z5895_assgn58956;
        z1951_assgn1951 <= z5895_assgn58957;
        z5901_assgn59010 <= z5901_assgn5901;
        z5901_assgn59011 <= z5901_assgn59010;
        z5901_assgn59012 <= z5901_assgn59011;
        z5901_assgn59013 <= z5901_assgn59012;
        z5901_assgn59014 <= z5901_assgn59013;
        z5901_assgn59015 <= z5901_assgn59014;
        z5901_assgn59016 <= z5901_assgn59015;
        z5901_assgn59017 <= z5901_assgn59016;
        z1955_assgn1955 <= z5901_assgn59017;
        z5939_assgn59390 <= z5939_assgn5939;
        z5939_assgn59391 <= z5939_assgn59390;
        z5939_assgn59392 <= z5939_assgn59391;
        z5939_assgn59393 <= z5939_assgn59392;
        z5939_assgn59394 <= z5939_assgn59393;
        z5939_assgn59395 <= z5939_assgn59394;
        z5939_assgn59396 <= z5939_assgn59395;
        z5939_assgn59397 <= z5939_assgn59396;
        z1991_assgn1991 <= z5939_assgn59397;
        z5945_assgn59450 <= z5945_assgn5945;
        z5945_assgn59451 <= z5945_assgn59450;
        z5945_assgn59452 <= z5945_assgn59451;
        z5945_assgn59453 <= z5945_assgn59452;
        z5945_assgn59454 <= z5945_assgn59453;
        z5945_assgn59455 <= z5945_assgn59454;
        z5945_assgn59456 <= z5945_assgn59455;
        z5945_assgn59457 <= z5945_assgn59456;
        z1995_assgn1995 <= z5945_assgn59457;
        z5951_assgn59510 <= z5951_assgn5951;
        z5951_assgn59511 <= z5951_assgn59510;
        z5951_assgn59512 <= z5951_assgn59511;
        z5951_assgn59513 <= z5951_assgn59512;
        z5951_assgn59514 <= z5951_assgn59513;
        z5951_assgn59515 <= z5951_assgn59514;
        z5951_assgn59516 <= z5951_assgn59515;
        z5951_assgn59517 <= z5951_assgn59516;
        z1999_assgn1999 <= z5951_assgn59517;
        z5993_assgn59930 <= z5993_assgn5993;
        z5993_assgn59931 <= z5993_assgn59930;
        z5993_assgn59932 <= z5993_assgn59931;
        z5993_assgn59933 <= z5993_assgn59932;
        z5993_assgn59934 <= z5993_assgn59933;
        z5993_assgn59935 <= z5993_assgn59934;
        z5993_assgn59936 <= z5993_assgn59935;
        z5993_assgn59937 <= z5993_assgn59936;
        z2039_assgn2039 <= z5993_assgn59937;
        m0_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= m0_comar0_G4_mul0_G16_mul1_G256_inv0;
        m1_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= m1_comar0_G4_mul0_G16_mul1_G256_inv0;
        z5999_assgn59990 <= z5999_assgn5999;
        z5999_assgn59991 <= z5999_assgn59990;
        z5999_assgn59992 <= z5999_assgn59991;
        z5999_assgn59993 <= z5999_assgn59992;
        z5999_assgn59994 <= z5999_assgn59993;
        z5999_assgn59995 <= z5999_assgn59994;
        z5999_assgn59996 <= z5999_assgn59995;
        z5999_assgn59997 <= z5999_assgn59996;
        z5999_assgn59998 <= z5999_assgn59997;
        z2043_assgn2043 <= z5999_assgn59998;
        m3_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= m3_comar0_G4_mul0_G16_mul1_G256_inv0;
        m2_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= m2_comar0_G4_mul0_G16_mul1_G256_inv0;
        z6005_assgn60050 <= z6005_assgn6005;
        z6005_assgn60051 <= z6005_assgn60050;
        z6005_assgn60052 <= z6005_assgn60051;
        z6005_assgn60053 <= z6005_assgn60052;
        z6005_assgn60054 <= z6005_assgn60053;
        z6005_assgn60055 <= z6005_assgn60054;
        z6005_assgn60056 <= z6005_assgn60055;
        z6005_assgn60057 <= z6005_assgn60056;
        z6005_assgn60058 <= z6005_assgn60057;
        z2047_assgn2047 <= z6005_assgn60058;
        r0_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= r0_10_comar0_G4_mul0_G16_mul1_G256_inv0;
        r1_10_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= r1_10_comar0_G4_mul0_G16_mul1_G256_inv0;
        z6013_assgn60130 <= z6013_assgn6013;
        z6013_assgn60131 <= z6013_assgn60130;
        z6013_assgn60132 <= z6013_assgn60131;
        z6013_assgn60133 <= z6013_assgn60132;
        z6013_assgn60134 <= z6013_assgn60133;
        z6013_assgn60135 <= z6013_assgn60134;
        z6013_assgn60136 <= z6013_assgn60135;
        z6013_assgn60137 <= z6013_assgn60136;
        z6013_assgn60138 <= z6013_assgn60137;
        z2053_assgn2053 <= z6013_assgn60138;
        z6017_assgn60170 <= z6017_assgn6017;
        z6017_assgn60171 <= z6017_assgn60170;
        z6017_assgn60172 <= z6017_assgn60171;
        z6017_assgn60173 <= z6017_assgn60172;
        z6017_assgn60174 <= z6017_assgn60173;
        z6017_assgn60175 <= z6017_assgn60174;
        z6017_assgn60176 <= z6017_assgn60175;
        z6017_assgn60177 <= z6017_assgn60176;
        z6017_assgn60178 <= z6017_assgn60177;
        z2055_assgn2055 <= z6017_assgn60178;
        z6021_assgn60210 <= z6021_assgn6021;
        z6021_assgn60211 <= z6021_assgn60210;
        z6021_assgn60212 <= z6021_assgn60211;
        z6021_assgn60213 <= z6021_assgn60212;
        z6021_assgn60214 <= z6021_assgn60213;
        z6021_assgn60215 <= z6021_assgn60214;
        z6021_assgn60216 <= z6021_assgn60215;
        z6021_assgn60217 <= z6021_assgn60216;
        z6021_assgn60218 <= z6021_assgn60217;
        z2058_assgn2058 <= z6021_assgn60218;
        i2_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= i2_comar0_G4_mul0_G16_mul1_G256_inv0;
        z6025_assgn60250 <= z6025_assgn6025;
        z6025_assgn60251 <= z6025_assgn60250;
        z6025_assgn60252 <= z6025_assgn60251;
        z6025_assgn60253 <= z6025_assgn60252;
        z6025_assgn60254 <= z6025_assgn60253;
        z6025_assgn60255 <= z6025_assgn60254;
        z6025_assgn60256 <= z6025_assgn60255;
        z6025_assgn60257 <= z6025_assgn60256;
        z6025_assgn60258 <= z6025_assgn60257;
        z2060_assgn2060 <= z6025_assgn60258;
        i3_comar0_G4_mul0_G16_mul1_G256_inv0_reg <= i3_comar0_G4_mul0_G16_mul1_G256_inv0;
        e0_G4_mul0_G16_mul1_G256_inv0 <= (i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0);
        z6059_assgn60590 <= z6059_assgn6059;
        z6059_assgn60591 <= z6059_assgn60590;
        z6059_assgn60592 <= z6059_assgn60591;
        z6059_assgn60593 <= z6059_assgn60592;
        z6059_assgn60594 <= z6059_assgn60593;
        z6059_assgn60595 <= z6059_assgn60594;
        z6059_assgn60596 <= z6059_assgn60595;
        z6059_assgn60597 <= z6059_assgn60596;
        z2091_assgn2091 <= z6059_assgn60597;
        m0_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= m0_comar1_G4_mul0_G16_mul1_G256_inv0;
        m1_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= m1_comar1_G4_mul0_G16_mul1_G256_inv0;
        z6065_assgn60650 <= z6065_assgn6065;
        z6065_assgn60651 <= z6065_assgn60650;
        z6065_assgn60652 <= z6065_assgn60651;
        z6065_assgn60653 <= z6065_assgn60652;
        z6065_assgn60654 <= z6065_assgn60653;
        z6065_assgn60655 <= z6065_assgn60654;
        z6065_assgn60656 <= z6065_assgn60655;
        z6065_assgn60657 <= z6065_assgn60656;
        z6065_assgn60658 <= z6065_assgn60657;
        z2095_assgn2095 <= z6065_assgn60658;
        m3_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= m3_comar1_G4_mul0_G16_mul1_G256_inv0;
        m2_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= m2_comar1_G4_mul0_G16_mul1_G256_inv0;
        z6071_assgn60710 <= z6071_assgn6071;
        z6071_assgn60711 <= z6071_assgn60710;
        z6071_assgn60712 <= z6071_assgn60711;
        z6071_assgn60713 <= z6071_assgn60712;
        z6071_assgn60714 <= z6071_assgn60713;
        z6071_assgn60715 <= z6071_assgn60714;
        z6071_assgn60716 <= z6071_assgn60715;
        z6071_assgn60717 <= z6071_assgn60716;
        z6071_assgn60718 <= z6071_assgn60717;
        z2099_assgn2099 <= z6071_assgn60718;
        r0_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= r0_10_comar1_G4_mul0_G16_mul1_G256_inv0;
        r1_10_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= r1_10_comar1_G4_mul0_G16_mul1_G256_inv0;
        z6079_assgn60790 <= z6079_assgn6079;
        z6079_assgn60791 <= z6079_assgn60790;
        z6079_assgn60792 <= z6079_assgn60791;
        z6079_assgn60793 <= z6079_assgn60792;
        z6079_assgn60794 <= z6079_assgn60793;
        z6079_assgn60795 <= z6079_assgn60794;
        z6079_assgn60796 <= z6079_assgn60795;
        z6079_assgn60797 <= z6079_assgn60796;
        z6079_assgn60798 <= z6079_assgn60797;
        z2105_assgn2105 <= z6079_assgn60798;
        z6083_assgn60830 <= z6083_assgn6083;
        z6083_assgn60831 <= z6083_assgn60830;
        z6083_assgn60832 <= z6083_assgn60831;
        z6083_assgn60833 <= z6083_assgn60832;
        z6083_assgn60834 <= z6083_assgn60833;
        z6083_assgn60835 <= z6083_assgn60834;
        z6083_assgn60836 <= z6083_assgn60835;
        z6083_assgn60837 <= z6083_assgn60836;
        z6083_assgn60838 <= z6083_assgn60837;
        z2107_assgn2107 <= z6083_assgn60838;
        z6087_assgn60870 <= z6087_assgn6087;
        z6087_assgn60871 <= z6087_assgn60870;
        z6087_assgn60872 <= z6087_assgn60871;
        z6087_assgn60873 <= z6087_assgn60872;
        z6087_assgn60874 <= z6087_assgn60873;
        z6087_assgn60875 <= z6087_assgn60874;
        z6087_assgn60876 <= z6087_assgn60875;
        z6087_assgn60877 <= z6087_assgn60876;
        z6087_assgn60878 <= z6087_assgn60877;
        z2110_assgn2110 <= z6087_assgn60878;
        i2_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= i2_comar1_G4_mul0_G16_mul1_G256_inv0;
        z6091_assgn60910 <= z6091_assgn6091;
        z6091_assgn60911 <= z6091_assgn60910;
        z6091_assgn60912 <= z6091_assgn60911;
        z6091_assgn60913 <= z6091_assgn60912;
        z6091_assgn60914 <= z6091_assgn60913;
        z6091_assgn60915 <= z6091_assgn60914;
        z6091_assgn60916 <= z6091_assgn60915;
        z6091_assgn60917 <= z6091_assgn60916;
        z6091_assgn60918 <= z6091_assgn60917;
        z2112_assgn2112 <= z6091_assgn60918;
        i3_comar1_G4_mul0_G16_mul1_G256_inv0_reg <= i3_comar1_G4_mul0_G16_mul1_G256_inv0;
        p0_0_G4_mul0_G16_mul1_G256_inv0 <= (i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0);
        z6129_assgn61290 <= z6129_assgn6129;
        z6129_assgn61291 <= z6129_assgn61290;
        z6129_assgn61292 <= z6129_assgn61291;
        z6129_assgn61293 <= z6129_assgn61292;
        z6129_assgn61294 <= z6129_assgn61293;
        z6129_assgn61295 <= z6129_assgn61294;
        z6129_assgn61296 <= z6129_assgn61295;
        z6129_assgn61297 <= z6129_assgn61296;
        z2147_assgn2147 <= z6129_assgn61297;
        m0_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= m0_comar2_G4_mul0_G16_mul1_G256_inv0;
        m1_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= m1_comar2_G4_mul0_G16_mul1_G256_inv0;
        z6135_assgn61350 <= z6135_assgn6135;
        z6135_assgn61351 <= z6135_assgn61350;
        z6135_assgn61352 <= z6135_assgn61351;
        z6135_assgn61353 <= z6135_assgn61352;
        z6135_assgn61354 <= z6135_assgn61353;
        z6135_assgn61355 <= z6135_assgn61354;
        z6135_assgn61356 <= z6135_assgn61355;
        z6135_assgn61357 <= z6135_assgn61356;
        z6135_assgn61358 <= z6135_assgn61357;
        z2151_assgn2151 <= z6135_assgn61358;
        m3_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= m3_comar2_G4_mul0_G16_mul1_G256_inv0;
        m2_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= m2_comar2_G4_mul0_G16_mul1_G256_inv0;
        z6141_assgn61410 <= z6141_assgn6141;
        z6141_assgn61411 <= z6141_assgn61410;
        z6141_assgn61412 <= z6141_assgn61411;
        z6141_assgn61413 <= z6141_assgn61412;
        z6141_assgn61414 <= z6141_assgn61413;
        z6141_assgn61415 <= z6141_assgn61414;
        z6141_assgn61416 <= z6141_assgn61415;
        z6141_assgn61417 <= z6141_assgn61416;
        z6141_assgn61418 <= z6141_assgn61417;
        z2155_assgn2155 <= z6141_assgn61418;
        r0_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= r0_10_comar2_G4_mul0_G16_mul1_G256_inv0;
        r1_10_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= r1_10_comar2_G4_mul0_G16_mul1_G256_inv0;
        z6149_assgn61490 <= z6149_assgn6149;
        z6149_assgn61491 <= z6149_assgn61490;
        z6149_assgn61492 <= z6149_assgn61491;
        z6149_assgn61493 <= z6149_assgn61492;
        z6149_assgn61494 <= z6149_assgn61493;
        z6149_assgn61495 <= z6149_assgn61494;
        z6149_assgn61496 <= z6149_assgn61495;
        z6149_assgn61497 <= z6149_assgn61496;
        z6149_assgn61498 <= z6149_assgn61497;
        z2161_assgn2161 <= z6149_assgn61498;
        z6153_assgn61530 <= z6153_assgn6153;
        z6153_assgn61531 <= z6153_assgn61530;
        z6153_assgn61532 <= z6153_assgn61531;
        z6153_assgn61533 <= z6153_assgn61532;
        z6153_assgn61534 <= z6153_assgn61533;
        z6153_assgn61535 <= z6153_assgn61534;
        z6153_assgn61536 <= z6153_assgn61535;
        z6153_assgn61537 <= z6153_assgn61536;
        z6153_assgn61538 <= z6153_assgn61537;
        z2163_assgn2163 <= z6153_assgn61538;
        z6157_assgn61570 <= z6157_assgn6157;
        z6157_assgn61571 <= z6157_assgn61570;
        z6157_assgn61572 <= z6157_assgn61571;
        z6157_assgn61573 <= z6157_assgn61572;
        z6157_assgn61574 <= z6157_assgn61573;
        z6157_assgn61575 <= z6157_assgn61574;
        z6157_assgn61576 <= z6157_assgn61575;
        z6157_assgn61577 <= z6157_assgn61576;
        z6157_assgn61578 <= z6157_assgn61577;
        z2166_assgn2166 <= z6157_assgn61578;
        i2_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= i2_comar2_G4_mul0_G16_mul1_G256_inv0;
        z6161_assgn61610 <= z6161_assgn6161;
        z6161_assgn61611 <= z6161_assgn61610;
        z6161_assgn61612 <= z6161_assgn61611;
        z6161_assgn61613 <= z6161_assgn61612;
        z6161_assgn61614 <= z6161_assgn61613;
        z6161_assgn61615 <= z6161_assgn61614;
        z6161_assgn61616 <= z6161_assgn61615;
        z6161_assgn61617 <= z6161_assgn61616;
        z6161_assgn61618 <= z6161_assgn61617;
        z2168_assgn2168 <= z6161_assgn61618;
        i3_comar2_G4_mul0_G16_mul1_G256_inv0_reg <= i3_comar2_G4_mul0_G16_mul1_G256_inv0;
        q0_0_G4_mul0_G16_mul1_G256_inv0 <= (i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0);
        z6183_assgn61830 <= z6183_assgn6183;
        z6183_assgn61831 <= z6183_assgn61830;
        z6183_assgn61832 <= z6183_assgn61831;
        z6183_assgn61833 <= z6183_assgn61832;
        z6183_assgn61834 <= z6183_assgn61833;
        z6183_assgn61835 <= z6183_assgn61834;
        z6183_assgn61836 <= z6183_assgn61835;
        z6183_assgn61837 <= z6183_assgn61836;
        z6183_assgn61838 <= z6183_assgn61837;
        z6183_assgn61839 <= z6183_assgn61838;
        z6183_assgn618310 <= z6183_assgn61839;
        z2187_assgn2187 <= z6183_assgn618310;
        z6193_assgn61930 <= z6193_assgn6193;
        z6193_assgn61931 <= z6193_assgn61930;
        z6193_assgn61932 <= z6193_assgn61931;
        z6193_assgn61933 <= z6193_assgn61932;
        z6193_assgn61934 <= z6193_assgn61933;
        z6193_assgn61935 <= z6193_assgn61934;
        z6193_assgn61936 <= z6193_assgn61935;
        z6193_assgn61937 <= z6193_assgn61936;
        z6193_assgn61938 <= z6193_assgn61937;
        z6193_assgn61939 <= z6193_assgn61938;
        z6193_assgn619310 <= z6193_assgn61939;
        z2195_assgn2195 <= z6193_assgn619310;
        z6199_assgn61990 <= z6199_assgn6199;
        z6199_assgn61991 <= z6199_assgn61990;
        z6199_assgn61992 <= z6199_assgn61991;
        z6199_assgn61993 <= z6199_assgn61992;
        z6199_assgn61994 <= z6199_assgn61993;
        z6199_assgn61995 <= z6199_assgn61994;
        z6199_assgn61996 <= z6199_assgn61995;
        z6199_assgn61997 <= z6199_assgn61996;
        z6199_assgn61998 <= z6199_assgn61997;
        z6199_assgn61999 <= z6199_assgn61998;
        z6199_assgn619910 <= z6199_assgn61999;
        z2199_assgn2199 <= z6199_assgn619910;
        z6205_assgn62050 <= z6205_assgn6205;
        z6205_assgn62051 <= z6205_assgn62050;
        z6205_assgn62052 <= z6205_assgn62051;
        z6205_assgn62053 <= z6205_assgn62052;
        z6205_assgn62054 <= z6205_assgn62053;
        z6205_assgn62055 <= z6205_assgn62054;
        z6205_assgn62056 <= z6205_assgn62055;
        z6205_assgn62057 <= z6205_assgn62056;
        z6205_assgn62058 <= z6205_assgn62057;
        z6205_assgn62059 <= z6205_assgn62058;
        z6205_assgn620510 <= z6205_assgn62059;
        z2203_assgn2203 <= z6205_assgn620510;
        z6217_assgn62170 <= z6217_assgn6217;
        z6217_assgn62171 <= z6217_assgn62170;
        z6217_assgn62172 <= z6217_assgn62171;
        z6217_assgn62173 <= z6217_assgn62172;
        z6217_assgn62174 <= z6217_assgn62173;
        z6217_assgn62175 <= z6217_assgn62174;
        z6217_assgn62176 <= z6217_assgn62175;
        z6217_assgn62177 <= z6217_assgn62176;
        z6217_assgn62178 <= z6217_assgn62177;
        z6217_assgn62179 <= z6217_assgn62178;
        z6217_assgn621710 <= z6217_assgn62179;
        z2213_assgn2213 <= z6217_assgn621710;
        z6241_assgn62410 <= z6241_assgn6241;
        z6241_assgn62411 <= z6241_assgn62410;
        z6241_assgn62412 <= z6241_assgn62411;
        z6241_assgn62413 <= z6241_assgn62412;
        z6241_assgn62414 <= z6241_assgn62413;
        z6241_assgn62415 <= z6241_assgn62414;
        z6241_assgn62416 <= z6241_assgn62415;
        z6241_assgn62417 <= z6241_assgn62416;
        z2235_assgn2235 <= z6241_assgn62417;
        z6247_assgn62470 <= z6247_assgn6247;
        z6247_assgn62471 <= z6247_assgn62470;
        z6247_assgn62472 <= z6247_assgn62471;
        z6247_assgn62473 <= z6247_assgn62472;
        z6247_assgn62474 <= z6247_assgn62473;
        z6247_assgn62475 <= z6247_assgn62474;
        z6247_assgn62476 <= z6247_assgn62475;
        z6247_assgn62477 <= z6247_assgn62476;
        z2239_assgn2239 <= z6247_assgn62477;
        z6253_assgn62530 <= z6253_assgn6253;
        z6253_assgn62531 <= z6253_assgn62530;
        z6253_assgn62532 <= z6253_assgn62531;
        z6253_assgn62533 <= z6253_assgn62532;
        z6253_assgn62534 <= z6253_assgn62533;
        z6253_assgn62535 <= z6253_assgn62534;
        z6253_assgn62536 <= z6253_assgn62535;
        z6253_assgn62537 <= z6253_assgn62536;
        z2243_assgn2243 <= z6253_assgn62537;
        z6295_assgn62950 <= z6295_assgn6295;
        z6295_assgn62951 <= z6295_assgn62950;
        z6295_assgn62952 <= z6295_assgn62951;
        z6295_assgn62953 <= z6295_assgn62952;
        z6295_assgn62954 <= z6295_assgn62953;
        z6295_assgn62955 <= z6295_assgn62954;
        z6295_assgn62956 <= z6295_assgn62955;
        z6295_assgn62957 <= z6295_assgn62956;
        z2283_assgn2283 <= z6295_assgn62957;
        m0_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= m0_comar0_G4_mul1_G16_mul1_G256_inv0;
        m1_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= m1_comar0_G4_mul1_G16_mul1_G256_inv0;
        z6301_assgn63010 <= z6301_assgn6301;
        z6301_assgn63011 <= z6301_assgn63010;
        z6301_assgn63012 <= z6301_assgn63011;
        z6301_assgn63013 <= z6301_assgn63012;
        z6301_assgn63014 <= z6301_assgn63013;
        z6301_assgn63015 <= z6301_assgn63014;
        z6301_assgn63016 <= z6301_assgn63015;
        z6301_assgn63017 <= z6301_assgn63016;
        z6301_assgn63018 <= z6301_assgn63017;
        z2287_assgn2287 <= z6301_assgn63018;
        m3_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= m3_comar0_G4_mul1_G16_mul1_G256_inv0;
        m2_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= m2_comar0_G4_mul1_G16_mul1_G256_inv0;
        z6307_assgn63070 <= z6307_assgn6307;
        z6307_assgn63071 <= z6307_assgn63070;
        z6307_assgn63072 <= z6307_assgn63071;
        z6307_assgn63073 <= z6307_assgn63072;
        z6307_assgn63074 <= z6307_assgn63073;
        z6307_assgn63075 <= z6307_assgn63074;
        z6307_assgn63076 <= z6307_assgn63075;
        z6307_assgn63077 <= z6307_assgn63076;
        z6307_assgn63078 <= z6307_assgn63077;
        z2291_assgn2291 <= z6307_assgn63078;
        r0_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= r0_10_comar0_G4_mul1_G16_mul1_G256_inv0;
        r1_10_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= r1_10_comar0_G4_mul1_G16_mul1_G256_inv0;
        z6315_assgn63150 <= z6315_assgn6315;
        z6315_assgn63151 <= z6315_assgn63150;
        z6315_assgn63152 <= z6315_assgn63151;
        z6315_assgn63153 <= z6315_assgn63152;
        z6315_assgn63154 <= z6315_assgn63153;
        z6315_assgn63155 <= z6315_assgn63154;
        z6315_assgn63156 <= z6315_assgn63155;
        z6315_assgn63157 <= z6315_assgn63156;
        z6315_assgn63158 <= z6315_assgn63157;
        z2297_assgn2297 <= z6315_assgn63158;
        z6319_assgn63190 <= z6319_assgn6319;
        z6319_assgn63191 <= z6319_assgn63190;
        z6319_assgn63192 <= z6319_assgn63191;
        z6319_assgn63193 <= z6319_assgn63192;
        z6319_assgn63194 <= z6319_assgn63193;
        z6319_assgn63195 <= z6319_assgn63194;
        z6319_assgn63196 <= z6319_assgn63195;
        z6319_assgn63197 <= z6319_assgn63196;
        z6319_assgn63198 <= z6319_assgn63197;
        z2299_assgn2299 <= z6319_assgn63198;
        z6323_assgn63230 <= z6323_assgn6323;
        z6323_assgn63231 <= z6323_assgn63230;
        z6323_assgn63232 <= z6323_assgn63231;
        z6323_assgn63233 <= z6323_assgn63232;
        z6323_assgn63234 <= z6323_assgn63233;
        z6323_assgn63235 <= z6323_assgn63234;
        z6323_assgn63236 <= z6323_assgn63235;
        z6323_assgn63237 <= z6323_assgn63236;
        z6323_assgn63238 <= z6323_assgn63237;
        z2302_assgn2302 <= z6323_assgn63238;
        i2_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= i2_comar0_G4_mul1_G16_mul1_G256_inv0;
        z6327_assgn63270 <= z6327_assgn6327;
        z6327_assgn63271 <= z6327_assgn63270;
        z6327_assgn63272 <= z6327_assgn63271;
        z6327_assgn63273 <= z6327_assgn63272;
        z6327_assgn63274 <= z6327_assgn63273;
        z6327_assgn63275 <= z6327_assgn63274;
        z6327_assgn63276 <= z6327_assgn63275;
        z6327_assgn63277 <= z6327_assgn63276;
        z6327_assgn63278 <= z6327_assgn63277;
        z2304_assgn2304 <= z6327_assgn63278;
        i3_comar0_G4_mul1_G16_mul1_G256_inv0_reg <= i3_comar0_G4_mul1_G16_mul1_G256_inv0;
        e0_G4_mul1_G16_mul1_G256_inv0 <= (i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0);
        z6361_assgn63610 <= z6361_assgn6361;
        z6361_assgn63611 <= z6361_assgn63610;
        z6361_assgn63612 <= z6361_assgn63611;
        z6361_assgn63613 <= z6361_assgn63612;
        z6361_assgn63614 <= z6361_assgn63613;
        z6361_assgn63615 <= z6361_assgn63614;
        z6361_assgn63616 <= z6361_assgn63615;
        z6361_assgn63617 <= z6361_assgn63616;
        z2335_assgn2335 <= z6361_assgn63617;
        m0_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= m0_comar1_G4_mul1_G16_mul1_G256_inv0;
        m1_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= m1_comar1_G4_mul1_G16_mul1_G256_inv0;
        z6367_assgn63670 <= z6367_assgn6367;
        z6367_assgn63671 <= z6367_assgn63670;
        z6367_assgn63672 <= z6367_assgn63671;
        z6367_assgn63673 <= z6367_assgn63672;
        z6367_assgn63674 <= z6367_assgn63673;
        z6367_assgn63675 <= z6367_assgn63674;
        z6367_assgn63676 <= z6367_assgn63675;
        z6367_assgn63677 <= z6367_assgn63676;
        z6367_assgn63678 <= z6367_assgn63677;
        z2339_assgn2339 <= z6367_assgn63678;
        m3_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= m3_comar1_G4_mul1_G16_mul1_G256_inv0;
        m2_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= m2_comar1_G4_mul1_G16_mul1_G256_inv0;
        z6373_assgn63730 <= z6373_assgn6373;
        z6373_assgn63731 <= z6373_assgn63730;
        z6373_assgn63732 <= z6373_assgn63731;
        z6373_assgn63733 <= z6373_assgn63732;
        z6373_assgn63734 <= z6373_assgn63733;
        z6373_assgn63735 <= z6373_assgn63734;
        z6373_assgn63736 <= z6373_assgn63735;
        z6373_assgn63737 <= z6373_assgn63736;
        z6373_assgn63738 <= z6373_assgn63737;
        z2343_assgn2343 <= z6373_assgn63738;
        r0_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= r0_10_comar1_G4_mul1_G16_mul1_G256_inv0;
        r1_10_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= r1_10_comar1_G4_mul1_G16_mul1_G256_inv0;
        z6381_assgn63810 <= z6381_assgn6381;
        z6381_assgn63811 <= z6381_assgn63810;
        z6381_assgn63812 <= z6381_assgn63811;
        z6381_assgn63813 <= z6381_assgn63812;
        z6381_assgn63814 <= z6381_assgn63813;
        z6381_assgn63815 <= z6381_assgn63814;
        z6381_assgn63816 <= z6381_assgn63815;
        z6381_assgn63817 <= z6381_assgn63816;
        z6381_assgn63818 <= z6381_assgn63817;
        z2349_assgn2349 <= z6381_assgn63818;
        z6385_assgn63850 <= z6385_assgn6385;
        z6385_assgn63851 <= z6385_assgn63850;
        z6385_assgn63852 <= z6385_assgn63851;
        z6385_assgn63853 <= z6385_assgn63852;
        z6385_assgn63854 <= z6385_assgn63853;
        z6385_assgn63855 <= z6385_assgn63854;
        z6385_assgn63856 <= z6385_assgn63855;
        z6385_assgn63857 <= z6385_assgn63856;
        z6385_assgn63858 <= z6385_assgn63857;
        z2351_assgn2351 <= z6385_assgn63858;
        z6389_assgn63890 <= z6389_assgn6389;
        z6389_assgn63891 <= z6389_assgn63890;
        z6389_assgn63892 <= z6389_assgn63891;
        z6389_assgn63893 <= z6389_assgn63892;
        z6389_assgn63894 <= z6389_assgn63893;
        z6389_assgn63895 <= z6389_assgn63894;
        z6389_assgn63896 <= z6389_assgn63895;
        z6389_assgn63897 <= z6389_assgn63896;
        z6389_assgn63898 <= z6389_assgn63897;
        z2354_assgn2354 <= z6389_assgn63898;
        i2_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= i2_comar1_G4_mul1_G16_mul1_G256_inv0;
        z6393_assgn63930 <= z6393_assgn6393;
        z6393_assgn63931 <= z6393_assgn63930;
        z6393_assgn63932 <= z6393_assgn63931;
        z6393_assgn63933 <= z6393_assgn63932;
        z6393_assgn63934 <= z6393_assgn63933;
        z6393_assgn63935 <= z6393_assgn63934;
        z6393_assgn63936 <= z6393_assgn63935;
        z6393_assgn63937 <= z6393_assgn63936;
        z6393_assgn63938 <= z6393_assgn63937;
        z2356_assgn2356 <= z6393_assgn63938;
        i3_comar1_G4_mul1_G16_mul1_G256_inv0_reg <= i3_comar1_G4_mul1_G16_mul1_G256_inv0;
        p0_0_G4_mul1_G16_mul1_G256_inv0 <= (i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0);
        z6431_assgn64310 <= z6431_assgn6431;
        z6431_assgn64311 <= z6431_assgn64310;
        z6431_assgn64312 <= z6431_assgn64311;
        z6431_assgn64313 <= z6431_assgn64312;
        z6431_assgn64314 <= z6431_assgn64313;
        z6431_assgn64315 <= z6431_assgn64314;
        z6431_assgn64316 <= z6431_assgn64315;
        z6431_assgn64317 <= z6431_assgn64316;
        z2391_assgn2391 <= z6431_assgn64317;
        m0_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= m0_comar2_G4_mul1_G16_mul1_G256_inv0;
        m1_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= m1_comar2_G4_mul1_G16_mul1_G256_inv0;
        z6437_assgn64370 <= z6437_assgn6437;
        z6437_assgn64371 <= z6437_assgn64370;
        z6437_assgn64372 <= z6437_assgn64371;
        z6437_assgn64373 <= z6437_assgn64372;
        z6437_assgn64374 <= z6437_assgn64373;
        z6437_assgn64375 <= z6437_assgn64374;
        z6437_assgn64376 <= z6437_assgn64375;
        z6437_assgn64377 <= z6437_assgn64376;
        z6437_assgn64378 <= z6437_assgn64377;
        z2395_assgn2395 <= z6437_assgn64378;
        m3_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= m3_comar2_G4_mul1_G16_mul1_G256_inv0;
        m2_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= m2_comar2_G4_mul1_G16_mul1_G256_inv0;
        z6443_assgn64430 <= z6443_assgn6443;
        z6443_assgn64431 <= z6443_assgn64430;
        z6443_assgn64432 <= z6443_assgn64431;
        z6443_assgn64433 <= z6443_assgn64432;
        z6443_assgn64434 <= z6443_assgn64433;
        z6443_assgn64435 <= z6443_assgn64434;
        z6443_assgn64436 <= z6443_assgn64435;
        z6443_assgn64437 <= z6443_assgn64436;
        z6443_assgn64438 <= z6443_assgn64437;
        z2399_assgn2399 <= z6443_assgn64438;
        r0_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= r0_10_comar2_G4_mul1_G16_mul1_G256_inv0;
        r1_10_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= r1_10_comar2_G4_mul1_G16_mul1_G256_inv0;
        z6451_assgn64510 <= z6451_assgn6451;
        z6451_assgn64511 <= z6451_assgn64510;
        z6451_assgn64512 <= z6451_assgn64511;
        z6451_assgn64513 <= z6451_assgn64512;
        z6451_assgn64514 <= z6451_assgn64513;
        z6451_assgn64515 <= z6451_assgn64514;
        z6451_assgn64516 <= z6451_assgn64515;
        z6451_assgn64517 <= z6451_assgn64516;
        z6451_assgn64518 <= z6451_assgn64517;
        z2405_assgn2405 <= z6451_assgn64518;
        z6455_assgn64550 <= z6455_assgn6455;
        z6455_assgn64551 <= z6455_assgn64550;
        z6455_assgn64552 <= z6455_assgn64551;
        z6455_assgn64553 <= z6455_assgn64552;
        z6455_assgn64554 <= z6455_assgn64553;
        z6455_assgn64555 <= z6455_assgn64554;
        z6455_assgn64556 <= z6455_assgn64555;
        z6455_assgn64557 <= z6455_assgn64556;
        z6455_assgn64558 <= z6455_assgn64557;
        z2407_assgn2407 <= z6455_assgn64558;
        z6459_assgn64590 <= z6459_assgn6459;
        z6459_assgn64591 <= z6459_assgn64590;
        z6459_assgn64592 <= z6459_assgn64591;
        z6459_assgn64593 <= z6459_assgn64592;
        z6459_assgn64594 <= z6459_assgn64593;
        z6459_assgn64595 <= z6459_assgn64594;
        z6459_assgn64596 <= z6459_assgn64595;
        z6459_assgn64597 <= z6459_assgn64596;
        z6459_assgn64598 <= z6459_assgn64597;
        z2410_assgn2410 <= z6459_assgn64598;
        i2_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= i2_comar2_G4_mul1_G16_mul1_G256_inv0;
        z6463_assgn64630 <= z6463_assgn6463;
        z6463_assgn64631 <= z6463_assgn64630;
        z6463_assgn64632 <= z6463_assgn64631;
        z6463_assgn64633 <= z6463_assgn64632;
        z6463_assgn64634 <= z6463_assgn64633;
        z6463_assgn64635 <= z6463_assgn64634;
        z6463_assgn64636 <= z6463_assgn64635;
        z6463_assgn64637 <= z6463_assgn64636;
        z6463_assgn64638 <= z6463_assgn64637;
        z2412_assgn2412 <= z6463_assgn64638;
        i3_comar2_G4_mul1_G16_mul1_G256_inv0_reg <= i3_comar2_G4_mul1_G16_mul1_G256_inv0;
        q0_0_G4_mul1_G16_mul1_G256_inv0 <= (i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0);
        z6485_assgn64850 <= z6485_assgn6485;
        z6485_assgn64851 <= z6485_assgn64850;
        z6485_assgn64852 <= z6485_assgn64851;
        z6485_assgn64853 <= z6485_assgn64852;
        z6485_assgn64854 <= z6485_assgn64853;
        z6485_assgn64855 <= z6485_assgn64854;
        z6485_assgn64856 <= z6485_assgn64855;
        z6485_assgn64857 <= z6485_assgn64856;
        z6485_assgn64858 <= z6485_assgn64857;
        z6485_assgn64859 <= z6485_assgn64858;
        z6485_assgn648510 <= z6485_assgn64859;
        z2431_assgn2431 <= z6485_assgn648510;
        z6511_assgn65110 <= z6511_assgn6511;
        z6511_assgn65111 <= z6511_assgn65110;
        z6511_assgn65112 <= z6511_assgn65111;
        z6511_assgn65113 <= z6511_assgn65112;
        z6511_assgn65114 <= z6511_assgn65113;
        z6511_assgn65115 <= z6511_assgn65114;
        z6511_assgn65116 <= z6511_assgn65115;
        z6511_assgn65117 <= z6511_assgn65116;
        z2455_assgn2455 <= z6511_assgn65117;
        z6517_assgn65170 <= z6517_assgn6517;
        z6517_assgn65171 <= z6517_assgn65170;
        z6517_assgn65172 <= z6517_assgn65171;
        z6517_assgn65173 <= z6517_assgn65172;
        z6517_assgn65174 <= z6517_assgn65173;
        z6517_assgn65175 <= z6517_assgn65174;
        z6517_assgn65176 <= z6517_assgn65175;
        z6517_assgn65177 <= z6517_assgn65176;
        z2459_assgn2459 <= z6517_assgn65177;
        z6523_assgn65230 <= z6523_assgn6523;
        z6523_assgn65231 <= z6523_assgn65230;
        z6523_assgn65232 <= z6523_assgn65231;
        z6523_assgn65233 <= z6523_assgn65232;
        z6523_assgn65234 <= z6523_assgn65233;
        z6523_assgn65235 <= z6523_assgn65234;
        z6523_assgn65236 <= z6523_assgn65235;
        z6523_assgn65237 <= z6523_assgn65236;
        z2463_assgn2463 <= z6523_assgn65237;
        z6565_assgn65650 <= z6565_assgn6565;
        z6565_assgn65651 <= z6565_assgn65650;
        z6565_assgn65652 <= z6565_assgn65651;
        z6565_assgn65653 <= z6565_assgn65652;
        z6565_assgn65654 <= z6565_assgn65653;
        z6565_assgn65655 <= z6565_assgn65654;
        z6565_assgn65656 <= z6565_assgn65655;
        z6565_assgn65657 <= z6565_assgn65656;
        z2503_assgn2503 <= z6565_assgn65657;
        m0_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= m0_comar0_G4_mul2_G16_mul1_G256_inv0;
        m1_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= m1_comar0_G4_mul2_G16_mul1_G256_inv0;
        z6571_assgn65710 <= z6571_assgn6571;
        z6571_assgn65711 <= z6571_assgn65710;
        z6571_assgn65712 <= z6571_assgn65711;
        z6571_assgn65713 <= z6571_assgn65712;
        z6571_assgn65714 <= z6571_assgn65713;
        z6571_assgn65715 <= z6571_assgn65714;
        z6571_assgn65716 <= z6571_assgn65715;
        z6571_assgn65717 <= z6571_assgn65716;
        z6571_assgn65718 <= z6571_assgn65717;
        z2507_assgn2507 <= z6571_assgn65718;
        m3_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= m3_comar0_G4_mul2_G16_mul1_G256_inv0;
        m2_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= m2_comar0_G4_mul2_G16_mul1_G256_inv0;
        z6577_assgn65770 <= z6577_assgn6577;
        z6577_assgn65771 <= z6577_assgn65770;
        z6577_assgn65772 <= z6577_assgn65771;
        z6577_assgn65773 <= z6577_assgn65772;
        z6577_assgn65774 <= z6577_assgn65773;
        z6577_assgn65775 <= z6577_assgn65774;
        z6577_assgn65776 <= z6577_assgn65775;
        z6577_assgn65777 <= z6577_assgn65776;
        z6577_assgn65778 <= z6577_assgn65777;
        z2511_assgn2511 <= z6577_assgn65778;
        r0_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= r0_10_comar0_G4_mul2_G16_mul1_G256_inv0;
        r1_10_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= r1_10_comar0_G4_mul2_G16_mul1_G256_inv0;
        z6585_assgn65850 <= z6585_assgn6585;
        z6585_assgn65851 <= z6585_assgn65850;
        z6585_assgn65852 <= z6585_assgn65851;
        z6585_assgn65853 <= z6585_assgn65852;
        z6585_assgn65854 <= z6585_assgn65853;
        z6585_assgn65855 <= z6585_assgn65854;
        z6585_assgn65856 <= z6585_assgn65855;
        z6585_assgn65857 <= z6585_assgn65856;
        z6585_assgn65858 <= z6585_assgn65857;
        z2517_assgn2517 <= z6585_assgn65858;
        z6589_assgn65890 <= z6589_assgn6589;
        z6589_assgn65891 <= z6589_assgn65890;
        z6589_assgn65892 <= z6589_assgn65891;
        z6589_assgn65893 <= z6589_assgn65892;
        z6589_assgn65894 <= z6589_assgn65893;
        z6589_assgn65895 <= z6589_assgn65894;
        z6589_assgn65896 <= z6589_assgn65895;
        z6589_assgn65897 <= z6589_assgn65896;
        z6589_assgn65898 <= z6589_assgn65897;
        z2519_assgn2519 <= z6589_assgn65898;
        z6593_assgn65930 <= z6593_assgn6593;
        z6593_assgn65931 <= z6593_assgn65930;
        z6593_assgn65932 <= z6593_assgn65931;
        z6593_assgn65933 <= z6593_assgn65932;
        z6593_assgn65934 <= z6593_assgn65933;
        z6593_assgn65935 <= z6593_assgn65934;
        z6593_assgn65936 <= z6593_assgn65935;
        z6593_assgn65937 <= z6593_assgn65936;
        z6593_assgn65938 <= z6593_assgn65937;
        z2522_assgn2522 <= z6593_assgn65938;
        i2_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= i2_comar0_G4_mul2_G16_mul1_G256_inv0;
        z6597_assgn65970 <= z6597_assgn6597;
        z6597_assgn65971 <= z6597_assgn65970;
        z6597_assgn65972 <= z6597_assgn65971;
        z6597_assgn65973 <= z6597_assgn65972;
        z6597_assgn65974 <= z6597_assgn65973;
        z6597_assgn65975 <= z6597_assgn65974;
        z6597_assgn65976 <= z6597_assgn65975;
        z6597_assgn65977 <= z6597_assgn65976;
        z6597_assgn65978 <= z6597_assgn65977;
        z2524_assgn2524 <= z6597_assgn65978;
        i3_comar0_G4_mul2_G16_mul1_G256_inv0_reg <= i3_comar0_G4_mul2_G16_mul1_G256_inv0;
        e0_G4_mul2_G16_mul1_G256_inv0 <= (i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0);
        z6631_assgn66310 <= z6631_assgn6631;
        z6631_assgn66311 <= z6631_assgn66310;
        z6631_assgn66312 <= z6631_assgn66311;
        z6631_assgn66313 <= z6631_assgn66312;
        z6631_assgn66314 <= z6631_assgn66313;
        z6631_assgn66315 <= z6631_assgn66314;
        z6631_assgn66316 <= z6631_assgn66315;
        z6631_assgn66317 <= z6631_assgn66316;
        z2555_assgn2555 <= z6631_assgn66317;
        m0_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= m0_comar1_G4_mul2_G16_mul1_G256_inv0;
        m1_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= m1_comar1_G4_mul2_G16_mul1_G256_inv0;
        z6637_assgn66370 <= z6637_assgn6637;
        z6637_assgn66371 <= z6637_assgn66370;
        z6637_assgn66372 <= z6637_assgn66371;
        z6637_assgn66373 <= z6637_assgn66372;
        z6637_assgn66374 <= z6637_assgn66373;
        z6637_assgn66375 <= z6637_assgn66374;
        z6637_assgn66376 <= z6637_assgn66375;
        z6637_assgn66377 <= z6637_assgn66376;
        z6637_assgn66378 <= z6637_assgn66377;
        z2559_assgn2559 <= z6637_assgn66378;
        m3_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= m3_comar1_G4_mul2_G16_mul1_G256_inv0;
        m2_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= m2_comar1_G4_mul2_G16_mul1_G256_inv0;
        z6643_assgn66430 <= z6643_assgn6643;
        z6643_assgn66431 <= z6643_assgn66430;
        z6643_assgn66432 <= z6643_assgn66431;
        z6643_assgn66433 <= z6643_assgn66432;
        z6643_assgn66434 <= z6643_assgn66433;
        z6643_assgn66435 <= z6643_assgn66434;
        z6643_assgn66436 <= z6643_assgn66435;
        z6643_assgn66437 <= z6643_assgn66436;
        z6643_assgn66438 <= z6643_assgn66437;
        z2563_assgn2563 <= z6643_assgn66438;
        r0_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= r0_10_comar1_G4_mul2_G16_mul1_G256_inv0;
        r1_10_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= r1_10_comar1_G4_mul2_G16_mul1_G256_inv0;
        z6651_assgn66510 <= z6651_assgn6651;
        z6651_assgn66511 <= z6651_assgn66510;
        z6651_assgn66512 <= z6651_assgn66511;
        z6651_assgn66513 <= z6651_assgn66512;
        z6651_assgn66514 <= z6651_assgn66513;
        z6651_assgn66515 <= z6651_assgn66514;
        z6651_assgn66516 <= z6651_assgn66515;
        z6651_assgn66517 <= z6651_assgn66516;
        z6651_assgn66518 <= z6651_assgn66517;
        z2569_assgn2569 <= z6651_assgn66518;
        z6655_assgn66550 <= z6655_assgn6655;
        z6655_assgn66551 <= z6655_assgn66550;
        z6655_assgn66552 <= z6655_assgn66551;
        z6655_assgn66553 <= z6655_assgn66552;
        z6655_assgn66554 <= z6655_assgn66553;
        z6655_assgn66555 <= z6655_assgn66554;
        z6655_assgn66556 <= z6655_assgn66555;
        z6655_assgn66557 <= z6655_assgn66556;
        z6655_assgn66558 <= z6655_assgn66557;
        z2571_assgn2571 <= z6655_assgn66558;
        z6659_assgn66590 <= z6659_assgn6659;
        z6659_assgn66591 <= z6659_assgn66590;
        z6659_assgn66592 <= z6659_assgn66591;
        z6659_assgn66593 <= z6659_assgn66592;
        z6659_assgn66594 <= z6659_assgn66593;
        z6659_assgn66595 <= z6659_assgn66594;
        z6659_assgn66596 <= z6659_assgn66595;
        z6659_assgn66597 <= z6659_assgn66596;
        z6659_assgn66598 <= z6659_assgn66597;
        z2574_assgn2574 <= z6659_assgn66598;
        i2_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= i2_comar1_G4_mul2_G16_mul1_G256_inv0;
        z6663_assgn66630 <= z6663_assgn6663;
        z6663_assgn66631 <= z6663_assgn66630;
        z6663_assgn66632 <= z6663_assgn66631;
        z6663_assgn66633 <= z6663_assgn66632;
        z6663_assgn66634 <= z6663_assgn66633;
        z6663_assgn66635 <= z6663_assgn66634;
        z6663_assgn66636 <= z6663_assgn66635;
        z6663_assgn66637 <= z6663_assgn66636;
        z6663_assgn66638 <= z6663_assgn66637;
        z2576_assgn2576 <= z6663_assgn66638;
        i3_comar1_G4_mul2_G16_mul1_G256_inv0_reg <= i3_comar1_G4_mul2_G16_mul1_G256_inv0;
        p0_0_G4_mul2_G16_mul1_G256_inv0 <= (i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0);
        z6701_assgn67010 <= z6701_assgn6701;
        z6701_assgn67011 <= z6701_assgn67010;
        z6701_assgn67012 <= z6701_assgn67011;
        z6701_assgn67013 <= z6701_assgn67012;
        z6701_assgn67014 <= z6701_assgn67013;
        z6701_assgn67015 <= z6701_assgn67014;
        z6701_assgn67016 <= z6701_assgn67015;
        z6701_assgn67017 <= z6701_assgn67016;
        z2611_assgn2611 <= z6701_assgn67017;
        m0_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= m0_comar2_G4_mul2_G16_mul1_G256_inv0;
        m1_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= m1_comar2_G4_mul2_G16_mul1_G256_inv0;
        z6707_assgn67070 <= z6707_assgn6707;
        z6707_assgn67071 <= z6707_assgn67070;
        z6707_assgn67072 <= z6707_assgn67071;
        z6707_assgn67073 <= z6707_assgn67072;
        z6707_assgn67074 <= z6707_assgn67073;
        z6707_assgn67075 <= z6707_assgn67074;
        z6707_assgn67076 <= z6707_assgn67075;
        z6707_assgn67077 <= z6707_assgn67076;
        z6707_assgn67078 <= z6707_assgn67077;
        z2615_assgn2615 <= z6707_assgn67078;
        m3_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= m3_comar2_G4_mul2_G16_mul1_G256_inv0;
        m2_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= m2_comar2_G4_mul2_G16_mul1_G256_inv0;
        z6713_assgn67130 <= z6713_assgn6713;
        z6713_assgn67131 <= z6713_assgn67130;
        z6713_assgn67132 <= z6713_assgn67131;
        z6713_assgn67133 <= z6713_assgn67132;
        z6713_assgn67134 <= z6713_assgn67133;
        z6713_assgn67135 <= z6713_assgn67134;
        z6713_assgn67136 <= z6713_assgn67135;
        z6713_assgn67137 <= z6713_assgn67136;
        z6713_assgn67138 <= z6713_assgn67137;
        z2619_assgn2619 <= z6713_assgn67138;
        r0_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= r0_10_comar2_G4_mul2_G16_mul1_G256_inv0;
        r1_10_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= r1_10_comar2_G4_mul2_G16_mul1_G256_inv0;
        z6721_assgn67210 <= z6721_assgn6721;
        z6721_assgn67211 <= z6721_assgn67210;
        z6721_assgn67212 <= z6721_assgn67211;
        z6721_assgn67213 <= z6721_assgn67212;
        z6721_assgn67214 <= z6721_assgn67213;
        z6721_assgn67215 <= z6721_assgn67214;
        z6721_assgn67216 <= z6721_assgn67215;
        z6721_assgn67217 <= z6721_assgn67216;
        z6721_assgn67218 <= z6721_assgn67217;
        z2625_assgn2625 <= z6721_assgn67218;
        z6725_assgn67250 <= z6725_assgn6725;
        z6725_assgn67251 <= z6725_assgn67250;
        z6725_assgn67252 <= z6725_assgn67251;
        z6725_assgn67253 <= z6725_assgn67252;
        z6725_assgn67254 <= z6725_assgn67253;
        z6725_assgn67255 <= z6725_assgn67254;
        z6725_assgn67256 <= z6725_assgn67255;
        z6725_assgn67257 <= z6725_assgn67256;
        z6725_assgn67258 <= z6725_assgn67257;
        z2627_assgn2627 <= z6725_assgn67258;
        z6729_assgn67290 <= z6729_assgn6729;
        z6729_assgn67291 <= z6729_assgn67290;
        z6729_assgn67292 <= z6729_assgn67291;
        z6729_assgn67293 <= z6729_assgn67292;
        z6729_assgn67294 <= z6729_assgn67293;
        z6729_assgn67295 <= z6729_assgn67294;
        z6729_assgn67296 <= z6729_assgn67295;
        z6729_assgn67297 <= z6729_assgn67296;
        z6729_assgn67298 <= z6729_assgn67297;
        z2630_assgn2630 <= z6729_assgn67298;
        i2_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= i2_comar2_G4_mul2_G16_mul1_G256_inv0;
        z6733_assgn67330 <= z6733_assgn6733;
        z6733_assgn67331 <= z6733_assgn67330;
        z6733_assgn67332 <= z6733_assgn67331;
        z6733_assgn67333 <= z6733_assgn67332;
        z6733_assgn67334 <= z6733_assgn67333;
        z6733_assgn67335 <= z6733_assgn67334;
        z6733_assgn67336 <= z6733_assgn67335;
        z6733_assgn67337 <= z6733_assgn67336;
        z6733_assgn67338 <= z6733_assgn67337;
        z2632_assgn2632 <= z6733_assgn67338;
        i3_comar2_G4_mul2_G16_mul1_G256_inv0_reg <= i3_comar2_G4_mul2_G16_mul1_G256_inv0;
        q0_0_G4_mul2_G16_mul1_G256_inv0 <= (i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0);
        z6755_assgn67550 <= z6755_assgn6755;
        z6755_assgn67551 <= z6755_assgn67550;
        z6755_assgn67552 <= z6755_assgn67551;
        z6755_assgn67553 <= z6755_assgn67552;
        z6755_assgn67554 <= z6755_assgn67553;
        z6755_assgn67555 <= z6755_assgn67554;
        z6755_assgn67556 <= z6755_assgn67555;
        z6755_assgn67557 <= z6755_assgn67556;
        z6755_assgn67558 <= z6755_assgn67557;
        z6755_assgn67559 <= z6755_assgn67558;
        z6755_assgn675510 <= z6755_assgn67559;
        z2651_assgn2651 <= z6755_assgn675510;
        z6769_assgn67690 <= z6769_assgn6769;
        z6769_assgn67691 <= z6769_assgn67690;
        z6769_assgn67692 <= z6769_assgn67691;
        z6769_assgn67693 <= z6769_assgn67692;
        z6769_assgn67694 <= z6769_assgn67693;
        z6769_assgn67695 <= z6769_assgn67694;
        z6769_assgn67696 <= z6769_assgn67695;
        z6769_assgn67697 <= z6769_assgn67696;
        z6769_assgn67698 <= z6769_assgn67697;
        z6769_assgn67699 <= z6769_assgn67698;
        z6769_assgn676910 <= z6769_assgn67699;
        z2663_assgn2663 <= z6769_assgn676910;
        z6791_assgn67910 <= z6791_assgn6791;
        z6791_assgn67911 <= z6791_assgn67910;
        z6791_assgn67912 <= z6791_assgn67911;
        z6791_assgn67913 <= z6791_assgn67912;
        z6791_assgn67914 <= z6791_assgn67913;
        z6791_assgn67915 <= z6791_assgn67914;
        z6791_assgn67916 <= z6791_assgn67915;
        z6791_assgn67917 <= z6791_assgn67916;
        z2683_assgn2683 <= z6791_assgn67917;
        z6797_assgn67970 <= z6797_assgn6797;
        z6797_assgn67971 <= z6797_assgn67970;
        z6797_assgn67972 <= z6797_assgn67971;
        z6797_assgn67973 <= z6797_assgn67972;
        z6797_assgn67974 <= z6797_assgn67973;
        z6797_assgn67975 <= z6797_assgn67974;
        z6797_assgn67976 <= z6797_assgn67975;
        z6797_assgn67977 <= z6797_assgn67976;
        z2687_assgn2687 <= z6797_assgn67977;
        z6803_assgn68030 <= z6803_assgn6803;
        z6803_assgn68031 <= z6803_assgn68030;
        z6803_assgn68032 <= z6803_assgn68031;
        z6803_assgn68033 <= z6803_assgn68032;
        z6803_assgn68034 <= z6803_assgn68033;
        z6803_assgn68035 <= z6803_assgn68034;
        z6803_assgn68036 <= z6803_assgn68035;
        z6803_assgn68037 <= z6803_assgn68036;
        z2691_assgn2691 <= z6803_assgn68037;
        z6841_assgn68410 <= z6841_assgn6841;
        z6841_assgn68411 <= z6841_assgn68410;
        z6841_assgn68412 <= z6841_assgn68411;
        z6841_assgn68413 <= z6841_assgn68412;
        z6841_assgn68414 <= z6841_assgn68413;
        z6841_assgn68415 <= z6841_assgn68414;
        z6841_assgn68416 <= z6841_assgn68415;
        z6841_assgn68417 <= z6841_assgn68416;
        z2727_assgn2727 <= z6841_assgn68417;
        z6847_assgn68470 <= z6847_assgn6847;
        z6847_assgn68471 <= z6847_assgn68470;
        z6847_assgn68472 <= z6847_assgn68471;
        z6847_assgn68473 <= z6847_assgn68472;
        z6847_assgn68474 <= z6847_assgn68473;
        z6847_assgn68475 <= z6847_assgn68474;
        z6847_assgn68476 <= z6847_assgn68475;
        z6847_assgn68477 <= z6847_assgn68476;
        z2731_assgn2731 <= z6847_assgn68477;
        z6853_assgn68530 <= z6853_assgn6853;
        z6853_assgn68531 <= z6853_assgn68530;
        z6853_assgn68532 <= z6853_assgn68531;
        z6853_assgn68533 <= z6853_assgn68532;
        z6853_assgn68534 <= z6853_assgn68533;
        z6853_assgn68535 <= z6853_assgn68534;
        z6853_assgn68536 <= z6853_assgn68535;
        z6853_assgn68537 <= z6853_assgn68536;
        z2735_assgn2735 <= z6853_assgn68537;
        z6895_assgn68950 <= z6895_assgn6895;
        z6895_assgn68951 <= z6895_assgn68950;
        z6895_assgn68952 <= z6895_assgn68951;
        z6895_assgn68953 <= z6895_assgn68952;
        z6895_assgn68954 <= z6895_assgn68953;
        z6895_assgn68955 <= z6895_assgn68954;
        z6895_assgn68956 <= z6895_assgn68955;
        z6895_assgn68957 <= z6895_assgn68956;
        z2775_assgn2775 <= z6895_assgn68957;
        m0_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= m0_comar0_G4_mul0_G16_mul2_G256_inv0;
        m1_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= m1_comar0_G4_mul0_G16_mul2_G256_inv0;
        z6901_assgn69010 <= z6901_assgn6901;
        z6901_assgn69011 <= z6901_assgn69010;
        z6901_assgn69012 <= z6901_assgn69011;
        z6901_assgn69013 <= z6901_assgn69012;
        z6901_assgn69014 <= z6901_assgn69013;
        z6901_assgn69015 <= z6901_assgn69014;
        z6901_assgn69016 <= z6901_assgn69015;
        z6901_assgn69017 <= z6901_assgn69016;
        z6901_assgn69018 <= z6901_assgn69017;
        z2779_assgn2779 <= z6901_assgn69018;
        m3_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= m3_comar0_G4_mul0_G16_mul2_G256_inv0;
        m2_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= m2_comar0_G4_mul0_G16_mul2_G256_inv0;
        z6907_assgn69070 <= z6907_assgn6907;
        z6907_assgn69071 <= z6907_assgn69070;
        z6907_assgn69072 <= z6907_assgn69071;
        z6907_assgn69073 <= z6907_assgn69072;
        z6907_assgn69074 <= z6907_assgn69073;
        z6907_assgn69075 <= z6907_assgn69074;
        z6907_assgn69076 <= z6907_assgn69075;
        z6907_assgn69077 <= z6907_assgn69076;
        z6907_assgn69078 <= z6907_assgn69077;
        z2783_assgn2783 <= z6907_assgn69078;
        r0_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= r0_10_comar0_G4_mul0_G16_mul2_G256_inv0;
        r1_10_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= r1_10_comar0_G4_mul0_G16_mul2_G256_inv0;
        z6915_assgn69150 <= z6915_assgn6915;
        z6915_assgn69151 <= z6915_assgn69150;
        z6915_assgn69152 <= z6915_assgn69151;
        z6915_assgn69153 <= z6915_assgn69152;
        z6915_assgn69154 <= z6915_assgn69153;
        z6915_assgn69155 <= z6915_assgn69154;
        z6915_assgn69156 <= z6915_assgn69155;
        z6915_assgn69157 <= z6915_assgn69156;
        z6915_assgn69158 <= z6915_assgn69157;
        z2789_assgn2789 <= z6915_assgn69158;
        z6919_assgn69190 <= z6919_assgn6919;
        z6919_assgn69191 <= z6919_assgn69190;
        z6919_assgn69192 <= z6919_assgn69191;
        z6919_assgn69193 <= z6919_assgn69192;
        z6919_assgn69194 <= z6919_assgn69193;
        z6919_assgn69195 <= z6919_assgn69194;
        z6919_assgn69196 <= z6919_assgn69195;
        z6919_assgn69197 <= z6919_assgn69196;
        z6919_assgn69198 <= z6919_assgn69197;
        z2791_assgn2791 <= z6919_assgn69198;
        z6923_assgn69230 <= z6923_assgn6923;
        z6923_assgn69231 <= z6923_assgn69230;
        z6923_assgn69232 <= z6923_assgn69231;
        z6923_assgn69233 <= z6923_assgn69232;
        z6923_assgn69234 <= z6923_assgn69233;
        z6923_assgn69235 <= z6923_assgn69234;
        z6923_assgn69236 <= z6923_assgn69235;
        z6923_assgn69237 <= z6923_assgn69236;
        z6923_assgn69238 <= z6923_assgn69237;
        z2794_assgn2794 <= z6923_assgn69238;
        i2_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= i2_comar0_G4_mul0_G16_mul2_G256_inv0;
        z6927_assgn69270 <= z6927_assgn6927;
        z6927_assgn69271 <= z6927_assgn69270;
        z6927_assgn69272 <= z6927_assgn69271;
        z6927_assgn69273 <= z6927_assgn69272;
        z6927_assgn69274 <= z6927_assgn69273;
        z6927_assgn69275 <= z6927_assgn69274;
        z6927_assgn69276 <= z6927_assgn69275;
        z6927_assgn69277 <= z6927_assgn69276;
        z6927_assgn69278 <= z6927_assgn69277;
        z2796_assgn2796 <= z6927_assgn69278;
        i3_comar0_G4_mul0_G16_mul2_G256_inv0_reg <= i3_comar0_G4_mul0_G16_mul2_G256_inv0;
        e0_G4_mul0_G16_mul2_G256_inv0 <= (i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0);
        z6961_assgn69610 <= z6961_assgn6961;
        z6961_assgn69611 <= z6961_assgn69610;
        z6961_assgn69612 <= z6961_assgn69611;
        z6961_assgn69613 <= z6961_assgn69612;
        z6961_assgn69614 <= z6961_assgn69613;
        z6961_assgn69615 <= z6961_assgn69614;
        z6961_assgn69616 <= z6961_assgn69615;
        z6961_assgn69617 <= z6961_assgn69616;
        z2827_assgn2827 <= z6961_assgn69617;
        m0_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= m0_comar1_G4_mul0_G16_mul2_G256_inv0;
        m1_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= m1_comar1_G4_mul0_G16_mul2_G256_inv0;
        z6967_assgn69670 <= z6967_assgn6967;
        z6967_assgn69671 <= z6967_assgn69670;
        z6967_assgn69672 <= z6967_assgn69671;
        z6967_assgn69673 <= z6967_assgn69672;
        z6967_assgn69674 <= z6967_assgn69673;
        z6967_assgn69675 <= z6967_assgn69674;
        z6967_assgn69676 <= z6967_assgn69675;
        z6967_assgn69677 <= z6967_assgn69676;
        z6967_assgn69678 <= z6967_assgn69677;
        z2831_assgn2831 <= z6967_assgn69678;
        m3_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= m3_comar1_G4_mul0_G16_mul2_G256_inv0;
        m2_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= m2_comar1_G4_mul0_G16_mul2_G256_inv0;
        z6973_assgn69730 <= z6973_assgn6973;
        z6973_assgn69731 <= z6973_assgn69730;
        z6973_assgn69732 <= z6973_assgn69731;
        z6973_assgn69733 <= z6973_assgn69732;
        z6973_assgn69734 <= z6973_assgn69733;
        z6973_assgn69735 <= z6973_assgn69734;
        z6973_assgn69736 <= z6973_assgn69735;
        z6973_assgn69737 <= z6973_assgn69736;
        z6973_assgn69738 <= z6973_assgn69737;
        z2835_assgn2835 <= z6973_assgn69738;
        r0_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= r0_10_comar1_G4_mul0_G16_mul2_G256_inv0;
        r1_10_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= r1_10_comar1_G4_mul0_G16_mul2_G256_inv0;
        z6981_assgn69810 <= z6981_assgn6981;
        z6981_assgn69811 <= z6981_assgn69810;
        z6981_assgn69812 <= z6981_assgn69811;
        z6981_assgn69813 <= z6981_assgn69812;
        z6981_assgn69814 <= z6981_assgn69813;
        z6981_assgn69815 <= z6981_assgn69814;
        z6981_assgn69816 <= z6981_assgn69815;
        z6981_assgn69817 <= z6981_assgn69816;
        z6981_assgn69818 <= z6981_assgn69817;
        z2841_assgn2841 <= z6981_assgn69818;
        z6985_assgn69850 <= z6985_assgn6985;
        z6985_assgn69851 <= z6985_assgn69850;
        z6985_assgn69852 <= z6985_assgn69851;
        z6985_assgn69853 <= z6985_assgn69852;
        z6985_assgn69854 <= z6985_assgn69853;
        z6985_assgn69855 <= z6985_assgn69854;
        z6985_assgn69856 <= z6985_assgn69855;
        z6985_assgn69857 <= z6985_assgn69856;
        z6985_assgn69858 <= z6985_assgn69857;
        z2843_assgn2843 <= z6985_assgn69858;
        z6989_assgn69890 <= z6989_assgn6989;
        z6989_assgn69891 <= z6989_assgn69890;
        z6989_assgn69892 <= z6989_assgn69891;
        z6989_assgn69893 <= z6989_assgn69892;
        z6989_assgn69894 <= z6989_assgn69893;
        z6989_assgn69895 <= z6989_assgn69894;
        z6989_assgn69896 <= z6989_assgn69895;
        z6989_assgn69897 <= z6989_assgn69896;
        z6989_assgn69898 <= z6989_assgn69897;
        z2846_assgn2846 <= z6989_assgn69898;
        i2_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= i2_comar1_G4_mul0_G16_mul2_G256_inv0;
        z6993_assgn69930 <= z6993_assgn6993;
        z6993_assgn69931 <= z6993_assgn69930;
        z6993_assgn69932 <= z6993_assgn69931;
        z6993_assgn69933 <= z6993_assgn69932;
        z6993_assgn69934 <= z6993_assgn69933;
        z6993_assgn69935 <= z6993_assgn69934;
        z6993_assgn69936 <= z6993_assgn69935;
        z6993_assgn69937 <= z6993_assgn69936;
        z6993_assgn69938 <= z6993_assgn69937;
        z2848_assgn2848 <= z6993_assgn69938;
        i3_comar1_G4_mul0_G16_mul2_G256_inv0_reg <= i3_comar1_G4_mul0_G16_mul2_G256_inv0;
        p0_0_G4_mul0_G16_mul2_G256_inv0 <= (i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0);
        z7031_assgn70310 <= z7031_assgn7031;
        z7031_assgn70311 <= z7031_assgn70310;
        z7031_assgn70312 <= z7031_assgn70311;
        z7031_assgn70313 <= z7031_assgn70312;
        z7031_assgn70314 <= z7031_assgn70313;
        z7031_assgn70315 <= z7031_assgn70314;
        z7031_assgn70316 <= z7031_assgn70315;
        z7031_assgn70317 <= z7031_assgn70316;
        z2883_assgn2883 <= z7031_assgn70317;
        m0_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= m0_comar2_G4_mul0_G16_mul2_G256_inv0;
        m1_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= m1_comar2_G4_mul0_G16_mul2_G256_inv0;
        z7037_assgn70370 <= z7037_assgn7037;
        z7037_assgn70371 <= z7037_assgn70370;
        z7037_assgn70372 <= z7037_assgn70371;
        z7037_assgn70373 <= z7037_assgn70372;
        z7037_assgn70374 <= z7037_assgn70373;
        z7037_assgn70375 <= z7037_assgn70374;
        z7037_assgn70376 <= z7037_assgn70375;
        z7037_assgn70377 <= z7037_assgn70376;
        z7037_assgn70378 <= z7037_assgn70377;
        z2887_assgn2887 <= z7037_assgn70378;
        m3_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= m3_comar2_G4_mul0_G16_mul2_G256_inv0;
        m2_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= m2_comar2_G4_mul0_G16_mul2_G256_inv0;
        z7043_assgn70430 <= z7043_assgn7043;
        z7043_assgn70431 <= z7043_assgn70430;
        z7043_assgn70432 <= z7043_assgn70431;
        z7043_assgn70433 <= z7043_assgn70432;
        z7043_assgn70434 <= z7043_assgn70433;
        z7043_assgn70435 <= z7043_assgn70434;
        z7043_assgn70436 <= z7043_assgn70435;
        z7043_assgn70437 <= z7043_assgn70436;
        z7043_assgn70438 <= z7043_assgn70437;
        z2891_assgn2891 <= z7043_assgn70438;
        r0_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= r0_10_comar2_G4_mul0_G16_mul2_G256_inv0;
        r1_10_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= r1_10_comar2_G4_mul0_G16_mul2_G256_inv0;
        z7051_assgn70510 <= z7051_assgn7051;
        z7051_assgn70511 <= z7051_assgn70510;
        z7051_assgn70512 <= z7051_assgn70511;
        z7051_assgn70513 <= z7051_assgn70512;
        z7051_assgn70514 <= z7051_assgn70513;
        z7051_assgn70515 <= z7051_assgn70514;
        z7051_assgn70516 <= z7051_assgn70515;
        z7051_assgn70517 <= z7051_assgn70516;
        z7051_assgn70518 <= z7051_assgn70517;
        z2897_assgn2897 <= z7051_assgn70518;
        z7055_assgn70550 <= z7055_assgn7055;
        z7055_assgn70551 <= z7055_assgn70550;
        z7055_assgn70552 <= z7055_assgn70551;
        z7055_assgn70553 <= z7055_assgn70552;
        z7055_assgn70554 <= z7055_assgn70553;
        z7055_assgn70555 <= z7055_assgn70554;
        z7055_assgn70556 <= z7055_assgn70555;
        z7055_assgn70557 <= z7055_assgn70556;
        z7055_assgn70558 <= z7055_assgn70557;
        z2899_assgn2899 <= z7055_assgn70558;
        z7059_assgn70590 <= z7059_assgn7059;
        z7059_assgn70591 <= z7059_assgn70590;
        z7059_assgn70592 <= z7059_assgn70591;
        z7059_assgn70593 <= z7059_assgn70592;
        z7059_assgn70594 <= z7059_assgn70593;
        z7059_assgn70595 <= z7059_assgn70594;
        z7059_assgn70596 <= z7059_assgn70595;
        z7059_assgn70597 <= z7059_assgn70596;
        z7059_assgn70598 <= z7059_assgn70597;
        z2902_assgn2902 <= z7059_assgn70598;
        i2_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= i2_comar2_G4_mul0_G16_mul2_G256_inv0;
        z7063_assgn70630 <= z7063_assgn7063;
        z7063_assgn70631 <= z7063_assgn70630;
        z7063_assgn70632 <= z7063_assgn70631;
        z7063_assgn70633 <= z7063_assgn70632;
        z7063_assgn70634 <= z7063_assgn70633;
        z7063_assgn70635 <= z7063_assgn70634;
        z7063_assgn70636 <= z7063_assgn70635;
        z7063_assgn70637 <= z7063_assgn70636;
        z7063_assgn70638 <= z7063_assgn70637;
        z2904_assgn2904 <= z7063_assgn70638;
        i3_comar2_G4_mul0_G16_mul2_G256_inv0_reg <= i3_comar2_G4_mul0_G16_mul2_G256_inv0;
        q0_0_G4_mul0_G16_mul2_G256_inv0 <= (i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0);
        z7085_assgn70850 <= z7085_assgn7085;
        z7085_assgn70851 <= z7085_assgn70850;
        z7085_assgn70852 <= z7085_assgn70851;
        z7085_assgn70853 <= z7085_assgn70852;
        z7085_assgn70854 <= z7085_assgn70853;
        z7085_assgn70855 <= z7085_assgn70854;
        z7085_assgn70856 <= z7085_assgn70855;
        z7085_assgn70857 <= z7085_assgn70856;
        z7085_assgn70858 <= z7085_assgn70857;
        z7085_assgn70859 <= z7085_assgn70858;
        z7085_assgn708510 <= z7085_assgn70859;
        z2923_assgn2923 <= z7085_assgn708510;
        z7095_assgn70950 <= z7095_assgn7095;
        z7095_assgn70951 <= z7095_assgn70950;
        z7095_assgn70952 <= z7095_assgn70951;
        z7095_assgn70953 <= z7095_assgn70952;
        z7095_assgn70954 <= z7095_assgn70953;
        z7095_assgn70955 <= z7095_assgn70954;
        z7095_assgn70956 <= z7095_assgn70955;
        z7095_assgn70957 <= z7095_assgn70956;
        z7095_assgn70958 <= z7095_assgn70957;
        z7095_assgn70959 <= z7095_assgn70958;
        z7095_assgn709510 <= z7095_assgn70959;
        z2931_assgn2931 <= z7095_assgn709510;
        z7101_assgn71010 <= z7101_assgn7101;
        z7101_assgn71011 <= z7101_assgn71010;
        z7101_assgn71012 <= z7101_assgn71011;
        z7101_assgn71013 <= z7101_assgn71012;
        z7101_assgn71014 <= z7101_assgn71013;
        z7101_assgn71015 <= z7101_assgn71014;
        z7101_assgn71016 <= z7101_assgn71015;
        z7101_assgn71017 <= z7101_assgn71016;
        z7101_assgn71018 <= z7101_assgn71017;
        z7101_assgn71019 <= z7101_assgn71018;
        z7101_assgn710110 <= z7101_assgn71019;
        z2935_assgn2935 <= z7101_assgn710110;
        z7107_assgn71070 <= z7107_assgn7107;
        z7107_assgn71071 <= z7107_assgn71070;
        z7107_assgn71072 <= z7107_assgn71071;
        z7107_assgn71073 <= z7107_assgn71072;
        z7107_assgn71074 <= z7107_assgn71073;
        z7107_assgn71075 <= z7107_assgn71074;
        z7107_assgn71076 <= z7107_assgn71075;
        z7107_assgn71077 <= z7107_assgn71076;
        z7107_assgn71078 <= z7107_assgn71077;
        z7107_assgn71079 <= z7107_assgn71078;
        z7107_assgn710710 <= z7107_assgn71079;
        z2939_assgn2939 <= z7107_assgn710710;
        z7119_assgn71190 <= z7119_assgn7119;
        z7119_assgn71191 <= z7119_assgn71190;
        z7119_assgn71192 <= z7119_assgn71191;
        z7119_assgn71193 <= z7119_assgn71192;
        z7119_assgn71194 <= z7119_assgn71193;
        z7119_assgn71195 <= z7119_assgn71194;
        z7119_assgn71196 <= z7119_assgn71195;
        z7119_assgn71197 <= z7119_assgn71196;
        z7119_assgn71198 <= z7119_assgn71197;
        z7119_assgn71199 <= z7119_assgn71198;
        z7119_assgn711910 <= z7119_assgn71199;
        z2949_assgn2949 <= z7119_assgn711910;
        z7143_assgn71430 <= z7143_assgn7143;
        z7143_assgn71431 <= z7143_assgn71430;
        z7143_assgn71432 <= z7143_assgn71431;
        z7143_assgn71433 <= z7143_assgn71432;
        z7143_assgn71434 <= z7143_assgn71433;
        z7143_assgn71435 <= z7143_assgn71434;
        z7143_assgn71436 <= z7143_assgn71435;
        z7143_assgn71437 <= z7143_assgn71436;
        z2971_assgn2971 <= z7143_assgn71437;
        z7149_assgn71490 <= z7149_assgn7149;
        z7149_assgn71491 <= z7149_assgn71490;
        z7149_assgn71492 <= z7149_assgn71491;
        z7149_assgn71493 <= z7149_assgn71492;
        z7149_assgn71494 <= z7149_assgn71493;
        z7149_assgn71495 <= z7149_assgn71494;
        z7149_assgn71496 <= z7149_assgn71495;
        z7149_assgn71497 <= z7149_assgn71496;
        z2975_assgn2975 <= z7149_assgn71497;
        z7155_assgn71550 <= z7155_assgn7155;
        z7155_assgn71551 <= z7155_assgn71550;
        z7155_assgn71552 <= z7155_assgn71551;
        z7155_assgn71553 <= z7155_assgn71552;
        z7155_assgn71554 <= z7155_assgn71553;
        z7155_assgn71555 <= z7155_assgn71554;
        z7155_assgn71556 <= z7155_assgn71555;
        z7155_assgn71557 <= z7155_assgn71556;
        z2979_assgn2979 <= z7155_assgn71557;
        z7197_assgn71970 <= z7197_assgn7197;
        z7197_assgn71971 <= z7197_assgn71970;
        z7197_assgn71972 <= z7197_assgn71971;
        z7197_assgn71973 <= z7197_assgn71972;
        z7197_assgn71974 <= z7197_assgn71973;
        z7197_assgn71975 <= z7197_assgn71974;
        z7197_assgn71976 <= z7197_assgn71975;
        z7197_assgn71977 <= z7197_assgn71976;
        z3019_assgn3019 <= z7197_assgn71977;
        m0_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= m0_comar0_G4_mul1_G16_mul2_G256_inv0;
        m1_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= m1_comar0_G4_mul1_G16_mul2_G256_inv0;
        z7203_assgn72030 <= z7203_assgn7203;
        z7203_assgn72031 <= z7203_assgn72030;
        z7203_assgn72032 <= z7203_assgn72031;
        z7203_assgn72033 <= z7203_assgn72032;
        z7203_assgn72034 <= z7203_assgn72033;
        z7203_assgn72035 <= z7203_assgn72034;
        z7203_assgn72036 <= z7203_assgn72035;
        z7203_assgn72037 <= z7203_assgn72036;
        z7203_assgn72038 <= z7203_assgn72037;
        z3023_assgn3023 <= z7203_assgn72038;
        m3_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= m3_comar0_G4_mul1_G16_mul2_G256_inv0;
        m2_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= m2_comar0_G4_mul1_G16_mul2_G256_inv0;
        z7209_assgn72090 <= z7209_assgn7209;
        z7209_assgn72091 <= z7209_assgn72090;
        z7209_assgn72092 <= z7209_assgn72091;
        z7209_assgn72093 <= z7209_assgn72092;
        z7209_assgn72094 <= z7209_assgn72093;
        z7209_assgn72095 <= z7209_assgn72094;
        z7209_assgn72096 <= z7209_assgn72095;
        z7209_assgn72097 <= z7209_assgn72096;
        z7209_assgn72098 <= z7209_assgn72097;
        z3027_assgn3027 <= z7209_assgn72098;
        r0_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= r0_10_comar0_G4_mul1_G16_mul2_G256_inv0;
        r1_10_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= r1_10_comar0_G4_mul1_G16_mul2_G256_inv0;
        z7217_assgn72170 <= z7217_assgn7217;
        z7217_assgn72171 <= z7217_assgn72170;
        z7217_assgn72172 <= z7217_assgn72171;
        z7217_assgn72173 <= z7217_assgn72172;
        z7217_assgn72174 <= z7217_assgn72173;
        z7217_assgn72175 <= z7217_assgn72174;
        z7217_assgn72176 <= z7217_assgn72175;
        z7217_assgn72177 <= z7217_assgn72176;
        z7217_assgn72178 <= z7217_assgn72177;
        z3033_assgn3033 <= z7217_assgn72178;
        z7221_assgn72210 <= z7221_assgn7221;
        z7221_assgn72211 <= z7221_assgn72210;
        z7221_assgn72212 <= z7221_assgn72211;
        z7221_assgn72213 <= z7221_assgn72212;
        z7221_assgn72214 <= z7221_assgn72213;
        z7221_assgn72215 <= z7221_assgn72214;
        z7221_assgn72216 <= z7221_assgn72215;
        z7221_assgn72217 <= z7221_assgn72216;
        z7221_assgn72218 <= z7221_assgn72217;
        z3035_assgn3035 <= z7221_assgn72218;
        z7225_assgn72250 <= z7225_assgn7225;
        z7225_assgn72251 <= z7225_assgn72250;
        z7225_assgn72252 <= z7225_assgn72251;
        z7225_assgn72253 <= z7225_assgn72252;
        z7225_assgn72254 <= z7225_assgn72253;
        z7225_assgn72255 <= z7225_assgn72254;
        z7225_assgn72256 <= z7225_assgn72255;
        z7225_assgn72257 <= z7225_assgn72256;
        z7225_assgn72258 <= z7225_assgn72257;
        z3038_assgn3038 <= z7225_assgn72258;
        i2_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= i2_comar0_G4_mul1_G16_mul2_G256_inv0;
        z7229_assgn72290 <= z7229_assgn7229;
        z7229_assgn72291 <= z7229_assgn72290;
        z7229_assgn72292 <= z7229_assgn72291;
        z7229_assgn72293 <= z7229_assgn72292;
        z7229_assgn72294 <= z7229_assgn72293;
        z7229_assgn72295 <= z7229_assgn72294;
        z7229_assgn72296 <= z7229_assgn72295;
        z7229_assgn72297 <= z7229_assgn72296;
        z7229_assgn72298 <= z7229_assgn72297;
        z3040_assgn3040 <= z7229_assgn72298;
        i3_comar0_G4_mul1_G16_mul2_G256_inv0_reg <= i3_comar0_G4_mul1_G16_mul2_G256_inv0;
        e0_G4_mul1_G16_mul2_G256_inv0 <= (i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0);
        z7263_assgn72630 <= z7263_assgn7263;
        z7263_assgn72631 <= z7263_assgn72630;
        z7263_assgn72632 <= z7263_assgn72631;
        z7263_assgn72633 <= z7263_assgn72632;
        z7263_assgn72634 <= z7263_assgn72633;
        z7263_assgn72635 <= z7263_assgn72634;
        z7263_assgn72636 <= z7263_assgn72635;
        z7263_assgn72637 <= z7263_assgn72636;
        z3071_assgn3071 <= z7263_assgn72637;
        m0_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= m0_comar1_G4_mul1_G16_mul2_G256_inv0;
        m1_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= m1_comar1_G4_mul1_G16_mul2_G256_inv0;
        z7269_assgn72690 <= z7269_assgn7269;
        z7269_assgn72691 <= z7269_assgn72690;
        z7269_assgn72692 <= z7269_assgn72691;
        z7269_assgn72693 <= z7269_assgn72692;
        z7269_assgn72694 <= z7269_assgn72693;
        z7269_assgn72695 <= z7269_assgn72694;
        z7269_assgn72696 <= z7269_assgn72695;
        z7269_assgn72697 <= z7269_assgn72696;
        z7269_assgn72698 <= z7269_assgn72697;
        z3075_assgn3075 <= z7269_assgn72698;
        m3_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= m3_comar1_G4_mul1_G16_mul2_G256_inv0;
        m2_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= m2_comar1_G4_mul1_G16_mul2_G256_inv0;
        z7275_assgn72750 <= z7275_assgn7275;
        z7275_assgn72751 <= z7275_assgn72750;
        z7275_assgn72752 <= z7275_assgn72751;
        z7275_assgn72753 <= z7275_assgn72752;
        z7275_assgn72754 <= z7275_assgn72753;
        z7275_assgn72755 <= z7275_assgn72754;
        z7275_assgn72756 <= z7275_assgn72755;
        z7275_assgn72757 <= z7275_assgn72756;
        z7275_assgn72758 <= z7275_assgn72757;
        z3079_assgn3079 <= z7275_assgn72758;
        r0_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= r0_10_comar1_G4_mul1_G16_mul2_G256_inv0;
        r1_10_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= r1_10_comar1_G4_mul1_G16_mul2_G256_inv0;
        z7283_assgn72830 <= z7283_assgn7283;
        z7283_assgn72831 <= z7283_assgn72830;
        z7283_assgn72832 <= z7283_assgn72831;
        z7283_assgn72833 <= z7283_assgn72832;
        z7283_assgn72834 <= z7283_assgn72833;
        z7283_assgn72835 <= z7283_assgn72834;
        z7283_assgn72836 <= z7283_assgn72835;
        z7283_assgn72837 <= z7283_assgn72836;
        z7283_assgn72838 <= z7283_assgn72837;
        z3085_assgn3085 <= z7283_assgn72838;
        z7287_assgn72870 <= z7287_assgn7287;
        z7287_assgn72871 <= z7287_assgn72870;
        z7287_assgn72872 <= z7287_assgn72871;
        z7287_assgn72873 <= z7287_assgn72872;
        z7287_assgn72874 <= z7287_assgn72873;
        z7287_assgn72875 <= z7287_assgn72874;
        z7287_assgn72876 <= z7287_assgn72875;
        z7287_assgn72877 <= z7287_assgn72876;
        z7287_assgn72878 <= z7287_assgn72877;
        z3087_assgn3087 <= z7287_assgn72878;
        z7291_assgn72910 <= z7291_assgn7291;
        z7291_assgn72911 <= z7291_assgn72910;
        z7291_assgn72912 <= z7291_assgn72911;
        z7291_assgn72913 <= z7291_assgn72912;
        z7291_assgn72914 <= z7291_assgn72913;
        z7291_assgn72915 <= z7291_assgn72914;
        z7291_assgn72916 <= z7291_assgn72915;
        z7291_assgn72917 <= z7291_assgn72916;
        z7291_assgn72918 <= z7291_assgn72917;
        z3090_assgn3090 <= z7291_assgn72918;
        i2_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= i2_comar1_G4_mul1_G16_mul2_G256_inv0;
        z7295_assgn72950 <= z7295_assgn7295;
        z7295_assgn72951 <= z7295_assgn72950;
        z7295_assgn72952 <= z7295_assgn72951;
        z7295_assgn72953 <= z7295_assgn72952;
        z7295_assgn72954 <= z7295_assgn72953;
        z7295_assgn72955 <= z7295_assgn72954;
        z7295_assgn72956 <= z7295_assgn72955;
        z7295_assgn72957 <= z7295_assgn72956;
        z7295_assgn72958 <= z7295_assgn72957;
        z3092_assgn3092 <= z7295_assgn72958;
        i3_comar1_G4_mul1_G16_mul2_G256_inv0_reg <= i3_comar1_G4_mul1_G16_mul2_G256_inv0;
        p0_0_G4_mul1_G16_mul2_G256_inv0 <= (i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0);
        z7333_assgn73330 <= z7333_assgn7333;
        z7333_assgn73331 <= z7333_assgn73330;
        z7333_assgn73332 <= z7333_assgn73331;
        z7333_assgn73333 <= z7333_assgn73332;
        z7333_assgn73334 <= z7333_assgn73333;
        z7333_assgn73335 <= z7333_assgn73334;
        z7333_assgn73336 <= z7333_assgn73335;
        z7333_assgn73337 <= z7333_assgn73336;
        z3127_assgn3127 <= z7333_assgn73337;
        m0_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= m0_comar2_G4_mul1_G16_mul2_G256_inv0;
        m1_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= m1_comar2_G4_mul1_G16_mul2_G256_inv0;
        z7339_assgn73390 <= z7339_assgn7339;
        z7339_assgn73391 <= z7339_assgn73390;
        z7339_assgn73392 <= z7339_assgn73391;
        z7339_assgn73393 <= z7339_assgn73392;
        z7339_assgn73394 <= z7339_assgn73393;
        z7339_assgn73395 <= z7339_assgn73394;
        z7339_assgn73396 <= z7339_assgn73395;
        z7339_assgn73397 <= z7339_assgn73396;
        z7339_assgn73398 <= z7339_assgn73397;
        z3131_assgn3131 <= z7339_assgn73398;
        m3_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= m3_comar2_G4_mul1_G16_mul2_G256_inv0;
        m2_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= m2_comar2_G4_mul1_G16_mul2_G256_inv0;
        z7345_assgn73450 <= z7345_assgn7345;
        z7345_assgn73451 <= z7345_assgn73450;
        z7345_assgn73452 <= z7345_assgn73451;
        z7345_assgn73453 <= z7345_assgn73452;
        z7345_assgn73454 <= z7345_assgn73453;
        z7345_assgn73455 <= z7345_assgn73454;
        z7345_assgn73456 <= z7345_assgn73455;
        z7345_assgn73457 <= z7345_assgn73456;
        z7345_assgn73458 <= z7345_assgn73457;
        z3135_assgn3135 <= z7345_assgn73458;
        r0_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= r0_10_comar2_G4_mul1_G16_mul2_G256_inv0;
        r1_10_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= r1_10_comar2_G4_mul1_G16_mul2_G256_inv0;
        z7353_assgn73530 <= z7353_assgn7353;
        z7353_assgn73531 <= z7353_assgn73530;
        z7353_assgn73532 <= z7353_assgn73531;
        z7353_assgn73533 <= z7353_assgn73532;
        z7353_assgn73534 <= z7353_assgn73533;
        z7353_assgn73535 <= z7353_assgn73534;
        z7353_assgn73536 <= z7353_assgn73535;
        z7353_assgn73537 <= z7353_assgn73536;
        z7353_assgn73538 <= z7353_assgn73537;
        z3141_assgn3141 <= z7353_assgn73538;
        z7357_assgn73570 <= z7357_assgn7357;
        z7357_assgn73571 <= z7357_assgn73570;
        z7357_assgn73572 <= z7357_assgn73571;
        z7357_assgn73573 <= z7357_assgn73572;
        z7357_assgn73574 <= z7357_assgn73573;
        z7357_assgn73575 <= z7357_assgn73574;
        z7357_assgn73576 <= z7357_assgn73575;
        z7357_assgn73577 <= z7357_assgn73576;
        z7357_assgn73578 <= z7357_assgn73577;
        z3143_assgn3143 <= z7357_assgn73578;
        z7361_assgn73610 <= z7361_assgn7361;
        z7361_assgn73611 <= z7361_assgn73610;
        z7361_assgn73612 <= z7361_assgn73611;
        z7361_assgn73613 <= z7361_assgn73612;
        z7361_assgn73614 <= z7361_assgn73613;
        z7361_assgn73615 <= z7361_assgn73614;
        z7361_assgn73616 <= z7361_assgn73615;
        z7361_assgn73617 <= z7361_assgn73616;
        z7361_assgn73618 <= z7361_assgn73617;
        z3146_assgn3146 <= z7361_assgn73618;
        i2_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= i2_comar2_G4_mul1_G16_mul2_G256_inv0;
        z7365_assgn73650 <= z7365_assgn7365;
        z7365_assgn73651 <= z7365_assgn73650;
        z7365_assgn73652 <= z7365_assgn73651;
        z7365_assgn73653 <= z7365_assgn73652;
        z7365_assgn73654 <= z7365_assgn73653;
        z7365_assgn73655 <= z7365_assgn73654;
        z7365_assgn73656 <= z7365_assgn73655;
        z7365_assgn73657 <= z7365_assgn73656;
        z7365_assgn73658 <= z7365_assgn73657;
        z3148_assgn3148 <= z7365_assgn73658;
        i3_comar2_G4_mul1_G16_mul2_G256_inv0_reg <= i3_comar2_G4_mul1_G16_mul2_G256_inv0;
        q0_0_G4_mul1_G16_mul2_G256_inv0 <= (i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0);
        z7387_assgn73870 <= z7387_assgn7387;
        z7387_assgn73871 <= z7387_assgn73870;
        z7387_assgn73872 <= z7387_assgn73871;
        z7387_assgn73873 <= z7387_assgn73872;
        z7387_assgn73874 <= z7387_assgn73873;
        z7387_assgn73875 <= z7387_assgn73874;
        z7387_assgn73876 <= z7387_assgn73875;
        z7387_assgn73877 <= z7387_assgn73876;
        z7387_assgn73878 <= z7387_assgn73877;
        z7387_assgn73879 <= z7387_assgn73878;
        z7387_assgn738710 <= z7387_assgn73879;
        z3167_assgn3167 <= z7387_assgn738710;
        z7413_assgn74130 <= z7413_assgn7413;
        z7413_assgn74131 <= z7413_assgn74130;
        z7413_assgn74132 <= z7413_assgn74131;
        z7413_assgn74133 <= z7413_assgn74132;
        z7413_assgn74134 <= z7413_assgn74133;
        z7413_assgn74135 <= z7413_assgn74134;
        z7413_assgn74136 <= z7413_assgn74135;
        z7413_assgn74137 <= z7413_assgn74136;
        z3191_assgn3191 <= z7413_assgn74137;
        z7419_assgn74190 <= z7419_assgn7419;
        z7419_assgn74191 <= z7419_assgn74190;
        z7419_assgn74192 <= z7419_assgn74191;
        z7419_assgn74193 <= z7419_assgn74192;
        z7419_assgn74194 <= z7419_assgn74193;
        z7419_assgn74195 <= z7419_assgn74194;
        z7419_assgn74196 <= z7419_assgn74195;
        z7419_assgn74197 <= z7419_assgn74196;
        z3195_assgn3195 <= z7419_assgn74197;
        z7425_assgn74250 <= z7425_assgn7425;
        z7425_assgn74251 <= z7425_assgn74250;
        z7425_assgn74252 <= z7425_assgn74251;
        z7425_assgn74253 <= z7425_assgn74252;
        z7425_assgn74254 <= z7425_assgn74253;
        z7425_assgn74255 <= z7425_assgn74254;
        z7425_assgn74256 <= z7425_assgn74255;
        z7425_assgn74257 <= z7425_assgn74256;
        z3199_assgn3199 <= z7425_assgn74257;
        z7467_assgn74670 <= z7467_assgn7467;
        z7467_assgn74671 <= z7467_assgn74670;
        z7467_assgn74672 <= z7467_assgn74671;
        z7467_assgn74673 <= z7467_assgn74672;
        z7467_assgn74674 <= z7467_assgn74673;
        z7467_assgn74675 <= z7467_assgn74674;
        z7467_assgn74676 <= z7467_assgn74675;
        z7467_assgn74677 <= z7467_assgn74676;
        z3239_assgn3239 <= z7467_assgn74677;
        m0_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= m0_comar0_G4_mul2_G16_mul2_G256_inv0;
        m1_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= m1_comar0_G4_mul2_G16_mul2_G256_inv0;
        z7473_assgn74730 <= z7473_assgn7473;
        z7473_assgn74731 <= z7473_assgn74730;
        z7473_assgn74732 <= z7473_assgn74731;
        z7473_assgn74733 <= z7473_assgn74732;
        z7473_assgn74734 <= z7473_assgn74733;
        z7473_assgn74735 <= z7473_assgn74734;
        z7473_assgn74736 <= z7473_assgn74735;
        z7473_assgn74737 <= z7473_assgn74736;
        z7473_assgn74738 <= z7473_assgn74737;
        z3243_assgn3243 <= z7473_assgn74738;
        m3_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= m3_comar0_G4_mul2_G16_mul2_G256_inv0;
        m2_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= m2_comar0_G4_mul2_G16_mul2_G256_inv0;
        z7479_assgn74790 <= z7479_assgn7479;
        z7479_assgn74791 <= z7479_assgn74790;
        z7479_assgn74792 <= z7479_assgn74791;
        z7479_assgn74793 <= z7479_assgn74792;
        z7479_assgn74794 <= z7479_assgn74793;
        z7479_assgn74795 <= z7479_assgn74794;
        z7479_assgn74796 <= z7479_assgn74795;
        z7479_assgn74797 <= z7479_assgn74796;
        z7479_assgn74798 <= z7479_assgn74797;
        z3247_assgn3247 <= z7479_assgn74798;
        r0_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= r0_10_comar0_G4_mul2_G16_mul2_G256_inv0;
        r1_10_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= r1_10_comar0_G4_mul2_G16_mul2_G256_inv0;
        z7487_assgn74870 <= z7487_assgn7487;
        z7487_assgn74871 <= z7487_assgn74870;
        z7487_assgn74872 <= z7487_assgn74871;
        z7487_assgn74873 <= z7487_assgn74872;
        z7487_assgn74874 <= z7487_assgn74873;
        z7487_assgn74875 <= z7487_assgn74874;
        z7487_assgn74876 <= z7487_assgn74875;
        z7487_assgn74877 <= z7487_assgn74876;
        z7487_assgn74878 <= z7487_assgn74877;
        z3253_assgn3253 <= z7487_assgn74878;
        z7491_assgn74910 <= z7491_assgn7491;
        z7491_assgn74911 <= z7491_assgn74910;
        z7491_assgn74912 <= z7491_assgn74911;
        z7491_assgn74913 <= z7491_assgn74912;
        z7491_assgn74914 <= z7491_assgn74913;
        z7491_assgn74915 <= z7491_assgn74914;
        z7491_assgn74916 <= z7491_assgn74915;
        z7491_assgn74917 <= z7491_assgn74916;
        z7491_assgn74918 <= z7491_assgn74917;
        z3255_assgn3255 <= z7491_assgn74918;
        z7495_assgn74950 <= z7495_assgn7495;
        z7495_assgn74951 <= z7495_assgn74950;
        z7495_assgn74952 <= z7495_assgn74951;
        z7495_assgn74953 <= z7495_assgn74952;
        z7495_assgn74954 <= z7495_assgn74953;
        z7495_assgn74955 <= z7495_assgn74954;
        z7495_assgn74956 <= z7495_assgn74955;
        z7495_assgn74957 <= z7495_assgn74956;
        z7495_assgn74958 <= z7495_assgn74957;
        z3258_assgn3258 <= z7495_assgn74958;
        i2_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= i2_comar0_G4_mul2_G16_mul2_G256_inv0;
        z7499_assgn74990 <= z7499_assgn7499;
        z7499_assgn74991 <= z7499_assgn74990;
        z7499_assgn74992 <= z7499_assgn74991;
        z7499_assgn74993 <= z7499_assgn74992;
        z7499_assgn74994 <= z7499_assgn74993;
        z7499_assgn74995 <= z7499_assgn74994;
        z7499_assgn74996 <= z7499_assgn74995;
        z7499_assgn74997 <= z7499_assgn74996;
        z7499_assgn74998 <= z7499_assgn74997;
        z3260_assgn3260 <= z7499_assgn74998;
        i3_comar0_G4_mul2_G16_mul2_G256_inv0_reg <= i3_comar0_G4_mul2_G16_mul2_G256_inv0;
        e0_G4_mul2_G16_mul2_G256_inv0 <= (i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0);
        z7533_assgn75330 <= z7533_assgn7533;
        z7533_assgn75331 <= z7533_assgn75330;
        z7533_assgn75332 <= z7533_assgn75331;
        z7533_assgn75333 <= z7533_assgn75332;
        z7533_assgn75334 <= z7533_assgn75333;
        z7533_assgn75335 <= z7533_assgn75334;
        z7533_assgn75336 <= z7533_assgn75335;
        z7533_assgn75337 <= z7533_assgn75336;
        z3291_assgn3291 <= z7533_assgn75337;
        m0_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= m0_comar1_G4_mul2_G16_mul2_G256_inv0;
        m1_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= m1_comar1_G4_mul2_G16_mul2_G256_inv0;
        z7539_assgn75390 <= z7539_assgn7539;
        z7539_assgn75391 <= z7539_assgn75390;
        z7539_assgn75392 <= z7539_assgn75391;
        z7539_assgn75393 <= z7539_assgn75392;
        z7539_assgn75394 <= z7539_assgn75393;
        z7539_assgn75395 <= z7539_assgn75394;
        z7539_assgn75396 <= z7539_assgn75395;
        z7539_assgn75397 <= z7539_assgn75396;
        z7539_assgn75398 <= z7539_assgn75397;
        z3295_assgn3295 <= z7539_assgn75398;
        m3_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= m3_comar1_G4_mul2_G16_mul2_G256_inv0;
        m2_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= m2_comar1_G4_mul2_G16_mul2_G256_inv0;
        z7545_assgn75450 <= z7545_assgn7545;
        z7545_assgn75451 <= z7545_assgn75450;
        z7545_assgn75452 <= z7545_assgn75451;
        z7545_assgn75453 <= z7545_assgn75452;
        z7545_assgn75454 <= z7545_assgn75453;
        z7545_assgn75455 <= z7545_assgn75454;
        z7545_assgn75456 <= z7545_assgn75455;
        z7545_assgn75457 <= z7545_assgn75456;
        z7545_assgn75458 <= z7545_assgn75457;
        z3299_assgn3299 <= z7545_assgn75458;
        r0_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= r0_10_comar1_G4_mul2_G16_mul2_G256_inv0;
        r1_10_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= r1_10_comar1_G4_mul2_G16_mul2_G256_inv0;
        z7553_assgn75530 <= z7553_assgn7553;
        z7553_assgn75531 <= z7553_assgn75530;
        z7553_assgn75532 <= z7553_assgn75531;
        z7553_assgn75533 <= z7553_assgn75532;
        z7553_assgn75534 <= z7553_assgn75533;
        z7553_assgn75535 <= z7553_assgn75534;
        z7553_assgn75536 <= z7553_assgn75535;
        z7553_assgn75537 <= z7553_assgn75536;
        z7553_assgn75538 <= z7553_assgn75537;
        z3305_assgn3305 <= z7553_assgn75538;
        z7557_assgn75570 <= z7557_assgn7557;
        z7557_assgn75571 <= z7557_assgn75570;
        z7557_assgn75572 <= z7557_assgn75571;
        z7557_assgn75573 <= z7557_assgn75572;
        z7557_assgn75574 <= z7557_assgn75573;
        z7557_assgn75575 <= z7557_assgn75574;
        z7557_assgn75576 <= z7557_assgn75575;
        z7557_assgn75577 <= z7557_assgn75576;
        z7557_assgn75578 <= z7557_assgn75577;
        z3307_assgn3307 <= z7557_assgn75578;
        z7561_assgn75610 <= z7561_assgn7561;
        z7561_assgn75611 <= z7561_assgn75610;
        z7561_assgn75612 <= z7561_assgn75611;
        z7561_assgn75613 <= z7561_assgn75612;
        z7561_assgn75614 <= z7561_assgn75613;
        z7561_assgn75615 <= z7561_assgn75614;
        z7561_assgn75616 <= z7561_assgn75615;
        z7561_assgn75617 <= z7561_assgn75616;
        z7561_assgn75618 <= z7561_assgn75617;
        z3310_assgn3310 <= z7561_assgn75618;
        i2_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= i2_comar1_G4_mul2_G16_mul2_G256_inv0;
        z7565_assgn75650 <= z7565_assgn7565;
        z7565_assgn75651 <= z7565_assgn75650;
        z7565_assgn75652 <= z7565_assgn75651;
        z7565_assgn75653 <= z7565_assgn75652;
        z7565_assgn75654 <= z7565_assgn75653;
        z7565_assgn75655 <= z7565_assgn75654;
        z7565_assgn75656 <= z7565_assgn75655;
        z7565_assgn75657 <= z7565_assgn75656;
        z7565_assgn75658 <= z7565_assgn75657;
        z3312_assgn3312 <= z7565_assgn75658;
        i3_comar1_G4_mul2_G16_mul2_G256_inv0_reg <= i3_comar1_G4_mul2_G16_mul2_G256_inv0;
        p0_0_G4_mul2_G16_mul2_G256_inv0 <= (i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0);
        z7603_assgn76030 <= z7603_assgn7603;
        z7603_assgn76031 <= z7603_assgn76030;
        z7603_assgn76032 <= z7603_assgn76031;
        z7603_assgn76033 <= z7603_assgn76032;
        z7603_assgn76034 <= z7603_assgn76033;
        z7603_assgn76035 <= z7603_assgn76034;
        z7603_assgn76036 <= z7603_assgn76035;
        z7603_assgn76037 <= z7603_assgn76036;
        z3347_assgn3347 <= z7603_assgn76037;
        m0_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= m0_comar2_G4_mul2_G16_mul2_G256_inv0;
        m1_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= m1_comar2_G4_mul2_G16_mul2_G256_inv0;
        z7609_assgn76090 <= z7609_assgn7609;
        z7609_assgn76091 <= z7609_assgn76090;
        z7609_assgn76092 <= z7609_assgn76091;
        z7609_assgn76093 <= z7609_assgn76092;
        z7609_assgn76094 <= z7609_assgn76093;
        z7609_assgn76095 <= z7609_assgn76094;
        z7609_assgn76096 <= z7609_assgn76095;
        z7609_assgn76097 <= z7609_assgn76096;
        z7609_assgn76098 <= z7609_assgn76097;
        z3351_assgn3351 <= z7609_assgn76098;
        m3_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= m3_comar2_G4_mul2_G16_mul2_G256_inv0;
        m2_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= m2_comar2_G4_mul2_G16_mul2_G256_inv0;
        z7615_assgn76150 <= z7615_assgn7615;
        z7615_assgn76151 <= z7615_assgn76150;
        z7615_assgn76152 <= z7615_assgn76151;
        z7615_assgn76153 <= z7615_assgn76152;
        z7615_assgn76154 <= z7615_assgn76153;
        z7615_assgn76155 <= z7615_assgn76154;
        z7615_assgn76156 <= z7615_assgn76155;
        z7615_assgn76157 <= z7615_assgn76156;
        z7615_assgn76158 <= z7615_assgn76157;
        z3355_assgn3355 <= z7615_assgn76158;
        r0_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= r0_10_comar2_G4_mul2_G16_mul2_G256_inv0;
        r1_10_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= r1_10_comar2_G4_mul2_G16_mul2_G256_inv0;
        z7623_assgn76230 <= z7623_assgn7623;
        z7623_assgn76231 <= z7623_assgn76230;
        z7623_assgn76232 <= z7623_assgn76231;
        z7623_assgn76233 <= z7623_assgn76232;
        z7623_assgn76234 <= z7623_assgn76233;
        z7623_assgn76235 <= z7623_assgn76234;
        z7623_assgn76236 <= z7623_assgn76235;
        z7623_assgn76237 <= z7623_assgn76236;
        z7623_assgn76238 <= z7623_assgn76237;
        z3361_assgn3361 <= z7623_assgn76238;
        z7627_assgn76270 <= z7627_assgn7627;
        z7627_assgn76271 <= z7627_assgn76270;
        z7627_assgn76272 <= z7627_assgn76271;
        z7627_assgn76273 <= z7627_assgn76272;
        z7627_assgn76274 <= z7627_assgn76273;
        z7627_assgn76275 <= z7627_assgn76274;
        z7627_assgn76276 <= z7627_assgn76275;
        z7627_assgn76277 <= z7627_assgn76276;
        z7627_assgn76278 <= z7627_assgn76277;
        z3363_assgn3363 <= z7627_assgn76278;
        z7631_assgn76310 <= z7631_assgn7631;
        z7631_assgn76311 <= z7631_assgn76310;
        z7631_assgn76312 <= z7631_assgn76311;
        z7631_assgn76313 <= z7631_assgn76312;
        z7631_assgn76314 <= z7631_assgn76313;
        z7631_assgn76315 <= z7631_assgn76314;
        z7631_assgn76316 <= z7631_assgn76315;
        z7631_assgn76317 <= z7631_assgn76316;
        z7631_assgn76318 <= z7631_assgn76317;
        z3366_assgn3366 <= z7631_assgn76318;
        i2_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= i2_comar2_G4_mul2_G16_mul2_G256_inv0;
        z7635_assgn76350 <= z7635_assgn7635;
        z7635_assgn76351 <= z7635_assgn76350;
        z7635_assgn76352 <= z7635_assgn76351;
        z7635_assgn76353 <= z7635_assgn76352;
        z7635_assgn76354 <= z7635_assgn76353;
        z7635_assgn76355 <= z7635_assgn76354;
        z7635_assgn76356 <= z7635_assgn76355;
        z7635_assgn76357 <= z7635_assgn76356;
        z7635_assgn76358 <= z7635_assgn76357;
        z3368_assgn3368 <= z7635_assgn76358;
        i3_comar2_G4_mul2_G16_mul2_G256_inv0_reg <= i3_comar2_G4_mul2_G16_mul2_G256_inv0;
        q0_0_G4_mul2_G16_mul2_G256_inv0 <= (i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0);
        z7657_assgn76570 <= z7657_assgn7657;
        z7657_assgn76571 <= z7657_assgn76570;
        z7657_assgn76572 <= z7657_assgn76571;
        z7657_assgn76573 <= z7657_assgn76572;
        z7657_assgn76574 <= z7657_assgn76573;
        z7657_assgn76575 <= z7657_assgn76574;
        z7657_assgn76576 <= z7657_assgn76575;
        z7657_assgn76577 <= z7657_assgn76576;
        z7657_assgn76578 <= z7657_assgn76577;
        z7657_assgn76579 <= z7657_assgn76578;
        z7657_assgn765710 <= z7657_assgn76579;
        z3387_assgn3387 <= z7657_assgn765710;
        z7671_assgn76710 <= z7671_assgn7671;
        z7671_assgn76711 <= z7671_assgn76710;
        z7671_assgn76712 <= z7671_assgn76711;
        z7671_assgn76713 <= z7671_assgn76712;
        z7671_assgn76714 <= z7671_assgn76713;
        z7671_assgn76715 <= z7671_assgn76714;
        z7671_assgn76716 <= z7671_assgn76715;
        z7671_assgn76717 <= z7671_assgn76716;
        z7671_assgn76718 <= z7671_assgn76717;
        z7671_assgn76719 <= z7671_assgn76718;
        z7671_assgn767110 <= z7671_assgn76719;
        z3399_assgn3399 <= z7671_assgn767110;
        z7681_assgn76810 <= z7681_assgn7681;
        z7681_assgn76811 <= z7681_assgn76810;
        z7681_assgn76812 <= z7681_assgn76811;
        z7681_assgn76813 <= z7681_assgn76812;
        z7681_assgn76814 <= z7681_assgn76813;
        z7681_assgn76815 <= z7681_assgn76814;
        z7681_assgn76816 <= z7681_assgn76815;
        z7681_assgn76817 <= z7681_assgn76816;
        z7681_assgn76818 <= z7681_assgn76817;
        z7681_assgn76819 <= z7681_assgn76818;
        z7681_assgn768110 <= z7681_assgn76819;
        z3407_assgn3407 <= z7681_assgn768110;
        z7817_assgn78170 <= z7817_assgn7817;
        z7817_assgn78171 <= z7817_assgn78170;
        z7817_assgn78172 <= z7817_assgn78171;
        z7817_assgn78173 <= z7817_assgn78172;
        z7817_assgn78174 <= z7817_assgn78173;
        z7817_assgn78175 <= z7817_assgn78174;
        z7817_assgn78176 <= z7817_assgn78175;
        z7817_assgn78177 <= z7817_assgn78176;
        z7817_assgn78178 <= z7817_assgn78177;
        z7817_assgn78179 <= z7817_assgn78178;
        z7817_assgn781710 <= z7817_assgn78179;
        x8_G256_newbasis1 <= z7817_assgn781710;
        z7825_assgn78250 <= z7825_assgn7825;
        z7825_assgn78251 <= z7825_assgn78250;
        z7825_assgn78252 <= z7825_assgn78251;
        z7825_assgn78253 <= z7825_assgn78252;
        z7825_assgn78254 <= z7825_assgn78253;
        z7825_assgn78255 <= z7825_assgn78254;
        z7825_assgn78256 <= z7825_assgn78255;
        z7825_assgn78257 <= z7825_assgn78256;
        z7825_assgn78258 <= z7825_assgn78257;
        z7825_assgn78259 <= z7825_assgn78258;
        z7825_assgn782510 <= z7825_assgn78259;
        z3549_assgn3549 <= z7825_assgn782510;
        z7833_assgn78330 <= z7833_assgn7833;
        z7833_assgn78331 <= z7833_assgn78330;
        z7833_assgn78332 <= z7833_assgn78331;
        z7833_assgn78333 <= z7833_assgn78332;
        z7833_assgn78334 <= z7833_assgn78333;
        z7833_assgn78335 <= z7833_assgn78334;
        z7833_assgn78336 <= z7833_assgn78335;
        z7833_assgn78337 <= z7833_assgn78336;
        z7833_assgn78338 <= z7833_assgn78337;
        z7833_assgn78339 <= z7833_assgn78338;
        z7833_assgn783310 <= z7833_assgn78339;
        z3555_assgn3555 <= z7833_assgn783310;
        z7837_assgn78370 <= z7837_assgn7837;
        z7837_assgn78371 <= z7837_assgn78370;
        z7837_assgn78372 <= z7837_assgn78371;
        z7837_assgn78373 <= z7837_assgn78372;
        z7837_assgn78374 <= z7837_assgn78373;
        z7837_assgn78375 <= z7837_assgn78374;
        z7837_assgn78376 <= z7837_assgn78375;
        z7837_assgn78377 <= z7837_assgn78376;
        z7837_assgn78378 <= z7837_assgn78377;
        z7837_assgn78379 <= z7837_assgn78378;
        z7837_assgn783710 <= z7837_assgn78379;
        z3558_assgn3558 <= z7837_assgn783710;
        z7843_assgn78430 <= z7843_assgn7843;
        z7843_assgn78431 <= z7843_assgn78430;
        z7843_assgn78432 <= z7843_assgn78431;
        z7843_assgn78433 <= z7843_assgn78432;
        z7843_assgn78434 <= z7843_assgn78433;
        z7843_assgn78435 <= z7843_assgn78434;
        z7843_assgn78436 <= z7843_assgn78435;
        z7843_assgn78437 <= z7843_assgn78436;
        z7843_assgn78438 <= z7843_assgn78437;
        z7843_assgn78439 <= z7843_assgn78438;
        z7843_assgn784310 <= z7843_assgn78439;
        z3561_assgn3561 <= z7843_assgn784310;
        z7849_assgn78490 <= z7849_assgn7849;
        z7849_assgn78491 <= z7849_assgn78490;
        z7849_assgn78492 <= z7849_assgn78491;
        z7849_assgn78493 <= z7849_assgn78492;
        z7849_assgn78494 <= z7849_assgn78493;
        z7849_assgn78495 <= z7849_assgn78494;
        z7849_assgn78496 <= z7849_assgn78495;
        z7849_assgn78497 <= z7849_assgn78496;
        z7849_assgn78498 <= z7849_assgn78497;
        z7849_assgn78499 <= z7849_assgn78498;
        z7849_assgn784910 <= z7849_assgn78499;
        z3565_assgn3565 <= z7849_assgn784910;
        z7855_assgn78550 <= z7855_assgn7855;
        z7855_assgn78551 <= z7855_assgn78550;
        z7855_assgn78552 <= z7855_assgn78551;
        z7855_assgn78553 <= z7855_assgn78552;
        z7855_assgn78554 <= z7855_assgn78553;
        z7855_assgn78555 <= z7855_assgn78554;
        z7855_assgn78556 <= z7855_assgn78555;
        z7855_assgn78557 <= z7855_assgn78556;
        z7855_assgn78558 <= z7855_assgn78557;
        z7855_assgn78559 <= z7855_assgn78558;
        z7855_assgn785510 <= z7855_assgn78559;
        z3569_assgn3569 <= z7855_assgn785510;
        z7865_assgn78650 <= z7865_assgn7865;
        z7865_assgn78651 <= z7865_assgn78650;
        z7865_assgn78652 <= z7865_assgn78651;
        z7865_assgn78653 <= z7865_assgn78652;
        z7865_assgn78654 <= z7865_assgn78653;
        z7865_assgn78655 <= z7865_assgn78654;
        z7865_assgn78656 <= z7865_assgn78655;
        z7865_assgn78657 <= z7865_assgn78656;
        z7865_assgn78658 <= z7865_assgn78657;
        z7865_assgn78659 <= z7865_assgn78658;
        z7865_assgn786510 <= z7865_assgn78659;
        z3577_assgn3577 <= z7865_assgn786510;
        z7871_assgn78710 <= z7871_assgn7871;
        z7871_assgn78711 <= z7871_assgn78710;
        z7871_assgn78712 <= z7871_assgn78711;
        z7871_assgn78713 <= z7871_assgn78712;
        z7871_assgn78714 <= z7871_assgn78713;
        z7871_assgn78715 <= z7871_assgn78714;
        z7871_assgn78716 <= z7871_assgn78715;
        z7871_assgn78717 <= z7871_assgn78716;
        z7871_assgn78718 <= z7871_assgn78717;
        z7871_assgn78719 <= z7871_assgn78718;
        z7871_assgn787110 <= z7871_assgn78719;
        z3581_assgn3581 <= z7871_assgn787110;
        z7877_assgn78770 <= z7877_assgn7877;
        z7877_assgn78771 <= z7877_assgn78770;
        z7877_assgn78772 <= z7877_assgn78771;
        z7877_assgn78773 <= z7877_assgn78772;
        z7877_assgn78774 <= z7877_assgn78773;
        z7877_assgn78775 <= z7877_assgn78774;
        z7877_assgn78776 <= z7877_assgn78775;
        z7877_assgn78777 <= z7877_assgn78776;
        z7877_assgn78778 <= z7877_assgn78777;
        z7877_assgn78779 <= z7877_assgn78778;
        z7877_assgn787710 <= z7877_assgn78779;
        z3585_assgn3585 <= z7877_assgn787710;
        z7887_assgn78870 <= z7887_assgn7887;
        z7887_assgn78871 <= z7887_assgn78870;
        z7887_assgn78872 <= z7887_assgn78871;
        z7887_assgn78873 <= z7887_assgn78872;
        z7887_assgn78874 <= z7887_assgn78873;
        z7887_assgn78875 <= z7887_assgn78874;
        z7887_assgn78876 <= z7887_assgn78875;
        z7887_assgn78877 <= z7887_assgn78876;
        z7887_assgn78878 <= z7887_assgn78877;
        z7887_assgn78879 <= z7887_assgn78878;
        z7887_assgn788710 <= z7887_assgn78879;
        z3593_assgn3593 <= z7887_assgn788710;
        z7893_assgn78930 <= z7893_assgn7893;
        z7893_assgn78931 <= z7893_assgn78930;
        z7893_assgn78932 <= z7893_assgn78931;
        z7893_assgn78933 <= z7893_assgn78932;
        z7893_assgn78934 <= z7893_assgn78933;
        z7893_assgn78935 <= z7893_assgn78934;
        z7893_assgn78936 <= z7893_assgn78935;
        z7893_assgn78937 <= z7893_assgn78936;
        z7893_assgn78938 <= z7893_assgn78937;
        z7893_assgn78939 <= z7893_assgn78938;
        z7893_assgn789310 <= z7893_assgn78939;
        z3597_assgn3597 <= z7893_assgn789310;
        z7899_assgn78990 <= z7899_assgn7899;
        z7899_assgn78991 <= z7899_assgn78990;
        z7899_assgn78992 <= z7899_assgn78991;
        z7899_assgn78993 <= z7899_assgn78992;
        z7899_assgn78994 <= z7899_assgn78993;
        z7899_assgn78995 <= z7899_assgn78994;
        z7899_assgn78996 <= z7899_assgn78995;
        z7899_assgn78997 <= z7899_assgn78996;
        z7899_assgn78998 <= z7899_assgn78997;
        z7899_assgn78999 <= z7899_assgn78998;
        z7899_assgn789910 <= z7899_assgn78999;
        z3601_assgn3601 <= z7899_assgn789910;
        z7909_assgn79090 <= z7909_assgn7909;
        z7909_assgn79091 <= z7909_assgn79090;
        z7909_assgn79092 <= z7909_assgn79091;
        z7909_assgn79093 <= z7909_assgn79092;
        z7909_assgn79094 <= z7909_assgn79093;
        z7909_assgn79095 <= z7909_assgn79094;
        z7909_assgn79096 <= z7909_assgn79095;
        z7909_assgn79097 <= z7909_assgn79096;
        z7909_assgn79098 <= z7909_assgn79097;
        z7909_assgn79099 <= z7909_assgn79098;
        z7909_assgn790910 <= z7909_assgn79099;
        z3609_assgn3609 <= z7909_assgn790910;
        z7915_assgn79150 <= z7915_assgn7915;
        z7915_assgn79151 <= z7915_assgn79150;
        z7915_assgn79152 <= z7915_assgn79151;
        z7915_assgn79153 <= z7915_assgn79152;
        z7915_assgn79154 <= z7915_assgn79153;
        z7915_assgn79155 <= z7915_assgn79154;
        z7915_assgn79156 <= z7915_assgn79155;
        z7915_assgn79157 <= z7915_assgn79156;
        z7915_assgn79158 <= z7915_assgn79157;
        z7915_assgn79159 <= z7915_assgn79158;
        z7915_assgn791510 <= z7915_assgn79159;
        z3613_assgn3613 <= z7915_assgn791510;
        z7921_assgn79210 <= z7921_assgn7921;
        z7921_assgn79211 <= z7921_assgn79210;
        z7921_assgn79212 <= z7921_assgn79211;
        z7921_assgn79213 <= z7921_assgn79212;
        z7921_assgn79214 <= z7921_assgn79213;
        z7921_assgn79215 <= z7921_assgn79214;
        z7921_assgn79216 <= z7921_assgn79215;
        z7921_assgn79217 <= z7921_assgn79216;
        z7921_assgn79218 <= z7921_assgn79217;
        z7921_assgn79219 <= z7921_assgn79218;
        z7921_assgn792110 <= z7921_assgn79219;
        z3617_assgn3617 <= z7921_assgn792110;
        z7931_assgn79310 <= z7931_assgn7931;
        z7931_assgn79311 <= z7931_assgn79310;
        z7931_assgn79312 <= z7931_assgn79311;
        z7931_assgn79313 <= z7931_assgn79312;
        z7931_assgn79314 <= z7931_assgn79313;
        z7931_assgn79315 <= z7931_assgn79314;
        z7931_assgn79316 <= z7931_assgn79315;
        z7931_assgn79317 <= z7931_assgn79316;
        z7931_assgn79318 <= z7931_assgn79317;
        z7931_assgn79319 <= z7931_assgn79318;
        z7931_assgn793110 <= z7931_assgn79319;
        z3625_assgn3625 <= z7931_assgn793110;
        z7937_assgn79370 <= z7937_assgn7937;
        z7937_assgn79371 <= z7937_assgn79370;
        z7937_assgn79372 <= z7937_assgn79371;
        z7937_assgn79373 <= z7937_assgn79372;
        z7937_assgn79374 <= z7937_assgn79373;
        z7937_assgn79375 <= z7937_assgn79374;
        z7937_assgn79376 <= z7937_assgn79375;
        z7937_assgn79377 <= z7937_assgn79376;
        z7937_assgn79378 <= z7937_assgn79377;
        z7937_assgn79379 <= z7937_assgn79378;
        z7937_assgn793710 <= z7937_assgn79379;
        z3629_assgn3629 <= z7937_assgn793710;
        z7943_assgn79430 <= z7943_assgn7943;
        z7943_assgn79431 <= z7943_assgn79430;
        z7943_assgn79432 <= z7943_assgn79431;
        z7943_assgn79433 <= z7943_assgn79432;
        z7943_assgn79434 <= z7943_assgn79433;
        z7943_assgn79435 <= z7943_assgn79434;
        z7943_assgn79436 <= z7943_assgn79435;
        z7943_assgn79437 <= z7943_assgn79436;
        z7943_assgn79438 <= z7943_assgn79437;
        z7943_assgn79439 <= z7943_assgn79438;
        z7943_assgn794310 <= z7943_assgn79439;
        z3633_assgn3633 <= z7943_assgn794310;
        z7953_assgn79530 <= z7953_assgn7953;
        z7953_assgn79531 <= z7953_assgn79530;
        z7953_assgn79532 <= z7953_assgn79531;
        z7953_assgn79533 <= z7953_assgn79532;
        z7953_assgn79534 <= z7953_assgn79533;
        z7953_assgn79535 <= z7953_assgn79534;
        z7953_assgn79536 <= z7953_assgn79535;
        z7953_assgn79537 <= z7953_assgn79536;
        z7953_assgn79538 <= z7953_assgn79537;
        z7953_assgn79539 <= z7953_assgn79538;
        z7953_assgn795310 <= z7953_assgn79539;
        z3641_assgn3641 <= z7953_assgn795310;
        z7959_assgn79590 <= z7959_assgn7959;
        z7959_assgn79591 <= z7959_assgn79590;
        z7959_assgn79592 <= z7959_assgn79591;
        z7959_assgn79593 <= z7959_assgn79592;
        z7959_assgn79594 <= z7959_assgn79593;
        z7959_assgn79595 <= z7959_assgn79594;
        z7959_assgn79596 <= z7959_assgn79595;
        z7959_assgn79597 <= z7959_assgn79596;
        z7959_assgn79598 <= z7959_assgn79597;
        z7959_assgn79599 <= z7959_assgn79598;
        z7959_assgn795910 <= z7959_assgn79599;
        z3645_assgn3645 <= z7959_assgn795910;
        z7965_assgn79650 <= z7965_assgn7965;
        z7965_assgn79651 <= z7965_assgn79650;
        z7965_assgn79652 <= z7965_assgn79651;
        z7965_assgn79653 <= z7965_assgn79652;
        z7965_assgn79654 <= z7965_assgn79653;
        z7965_assgn79655 <= z7965_assgn79654;
        z7965_assgn79656 <= z7965_assgn79655;
        z7965_assgn79657 <= z7965_assgn79656;
        z7965_assgn79658 <= z7965_assgn79657;
        z7965_assgn79659 <= z7965_assgn79658;
        z7965_assgn796510 <= z7965_assgn79659;
        z3649_assgn3649 <= z7965_assgn796510;
        z7975_assgn79750 <= z7975_assgn7975;
        z7975_assgn79751 <= z7975_assgn79750;
        z7975_assgn79752 <= z7975_assgn79751;
        z7975_assgn79753 <= z7975_assgn79752;
        z7975_assgn79754 <= z7975_assgn79753;
        z7975_assgn79755 <= z7975_assgn79754;
        z7975_assgn79756 <= z7975_assgn79755;
        z7975_assgn79757 <= z7975_assgn79756;
        z7975_assgn79758 <= z7975_assgn79757;
        z7975_assgn79759 <= z7975_assgn79758;
        z7975_assgn797510 <= z7975_assgn79759;
        z3657_assgn3657 <= z7975_assgn797510;
        z7981_assgn79810 <= z7981_assgn7981;
        z7981_assgn79811 <= z7981_assgn79810;
        z7981_assgn79812 <= z7981_assgn79811;
        z7981_assgn79813 <= z7981_assgn79812;
        z7981_assgn79814 <= z7981_assgn79813;
        z7981_assgn79815 <= z7981_assgn79814;
        z7981_assgn79816 <= z7981_assgn79815;
        z7981_assgn79817 <= z7981_assgn79816;
        z7981_assgn79818 <= z7981_assgn79817;
        z7981_assgn79819 <= z7981_assgn79818;
        z7981_assgn798110 <= z7981_assgn79819;
        z3661_assgn3661 <= z7981_assgn798110;
        z7987_assgn79870 <= z7987_assgn7987;
        z7987_assgn79871 <= z7987_assgn79870;
        z7987_assgn79872 <= z7987_assgn79871;
        z7987_assgn79873 <= z7987_assgn79872;
        z7987_assgn79874 <= z7987_assgn79873;
        z7987_assgn79875 <= z7987_assgn79874;
        z7987_assgn79876 <= z7987_assgn79875;
        z7987_assgn79877 <= z7987_assgn79876;
        z7987_assgn79878 <= z7987_assgn79877;
        z7987_assgn79879 <= z7987_assgn79878;
        z7987_assgn798710 <= z7987_assgn79879;
        z3665_assgn3665 <= z7987_assgn798710;
        z7997_assgn79970 <= z7997_assgn7997;
        z7997_assgn79971 <= z7997_assgn79970;
        z7997_assgn79972 <= z7997_assgn79971;
        z7997_assgn79973 <= z7997_assgn79972;
        z7997_assgn79974 <= z7997_assgn79973;
        z7997_assgn79975 <= z7997_assgn79974;
        z7997_assgn79976 <= z7997_assgn79975;
        z7997_assgn79977 <= z7997_assgn79976;
        z7997_assgn79978 <= z7997_assgn79977;
        z7997_assgn79979 <= z7997_assgn79978;
        z7997_assgn799710 <= z7997_assgn79979;
        z3673_assgn3673 <= z7997_assgn799710;
        z8003_assgn80030 <= z8003_assgn8003;
        z8003_assgn80031 <= z8003_assgn80030;
        z8003_assgn80032 <= z8003_assgn80031;
        z8003_assgn80033 <= z8003_assgn80032;
        z8003_assgn80034 <= z8003_assgn80033;
        z8003_assgn80035 <= z8003_assgn80034;
        z8003_assgn80036 <= z8003_assgn80035;
        z8003_assgn80037 <= z8003_assgn80036;
        z8003_assgn80038 <= z8003_assgn80037;
        z8003_assgn80039 <= z8003_assgn80038;
        z8003_assgn800310 <= z8003_assgn80039;
        y0 <= z8003_assgn800310;
        y1 <= t7;
    end

endmodule

