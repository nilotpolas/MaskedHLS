module sbox(
    clk,
    x0_0,
    x1_0,
    x2_0,
    x3_0,
    x0_1,
    x1_1,
    x2_1,
    x3_1,
    r,
    Y0_0,
    Y1_0,
    Y2_0,
    Y3_0,
    Y0_1,
    Y1_1,
    Y2_1,
    Y3_1
);
//INPUTS
    input clk;
    input  x0_0;
    input  x1_0;
    input  x2_0;
    input  x3_0;
    input  x0_1;
    input  x1_1;
    input  x2_1;
    input  x3_1;
    input  r;
//OUTPUTS
    output reg  Y0_0;
    output reg  Y1_0;
    output reg  Y2_0;
    output reg  Y3_0;
    output reg  Y0_1;
    output reg  Y1_1;
    output reg  Y2_1;
    output reg  Y3_1;
//Intermediate values
    wire x0_0_inp;
    wire x1_0_inp;
    wire x2_0_inp;
    wire x3_0_inp;
    wire x0_1_inp;
    wire x1_1_inp;
    wire x2_1_inp;
    wire x3_1_inp;
    wire r_inp;
    wire L0_0;
    wire L1_0;
    wire L8_0;
    wire L5_0;
    wire L0_1;
    wire L1_1;
    wire L8_1;
    wire L5_1;
    wire Q0_0;
    wire Q1_0;
    wire Q3_0;
    wire Q4_0;
    wire Q0_1;
    wire Q1_1;
    wire Q3_1;
    wire Q4_1;
    wire L2_0;
    wire L3_0;
    wire L2_1;
    wire L3_1;
    wire p2_domand0;
    wire i1_domand0;
    wire p3_domand0;
    wire i2_domand0;
    wire p1_domand0;
    wire p4_domand0;
    reg i1_domand0_reg;
    reg p1_domand0_reg;
    wire T0_0;
    reg i2_domand0_reg;
    reg p4_domand0_reg;
    wire T0_1;
    wire L10_0;
    wire L10_1;
    wire p2_domand1;
    wire i1_domand1;
    wire p3_domand1;
    wire i2_domand1;
    wire p1_domand1;
    wire p4_domand1;
    reg i1_domand1_reg;
    reg p1_domand1_reg;
    wire T2_0;
    reg i2_domand1_reg;
    reg p4_domand1_reg;
    wire T2_1;
    reg L2_0_reg;
    wire Q2_0;
    wire L4_0;
    reg L5_0_reg;
    wire Q7_0;
    reg L3_0_reg;
    wire Q6_0;
    reg L2_1_reg;
    wire Q2_1;
    wire L4_1;
    reg L5_1_reg;
    wire Q7_1;
    reg L3_1_reg;
    wire Q6_1;
    reg Q3_1_reg;
    wire p2_domand2;
    reg r_inp_reg;
    wire i1_domand2;
    reg Q3_0_reg;
    wire p3_domand2;
    wire i2_domand2;
    wire p1_domand2;
    wire p4_domand2;
    reg i1_domand2_reg;
    reg p1_domand2_reg;
    wire T1_0;
    reg i2_domand2_reg;
    reg p4_domand2_reg;
    wire T1_1;
    wire p2_domand3;
    wire i1_domand3;
    wire p3_domand3;
    wire i2_domand3;
    wire p1_domand3;
    wire p4_domand3;
    reg i1_domand3_reg;
    reg p1_domand3_reg;
    wire T3_0;
    reg i2_domand3_reg;
    reg p4_domand3_reg;
    wire T3_1;
    reg T0_0_reg;
    wire L7_0;
    wire z343_assgn343;
    reg z343_assgn3430;
    reg z157_assgn157;
    wire L11_0;
    reg T0_1_reg;
    wire L7_1;
    wire z349_assgn349;
    reg z349_assgn3490;
    reg z161_assgn161;
    wire L11_1;
    reg T2_0_reg;
    wire Y0_01;
    wire z355_assgn355;
    reg z355_assgn3550;
    reg z166_assgn166;
    wire Y1_01;
    reg T2_1_reg;
    wire Y0_11;
    wire z361_assgn361;
    reg z361_assgn3610;
    reg z170_assgn170;
    wire Y1_11;
    wire z365_assgn365;
    reg z365_assgn3650;
    reg z172_assgn172;
    wire z1_assgn1;
    wire z3_assgn3;
    wire z5_assgn5;
    wire z379_assgn379;
    reg z379_assgn3790;
    wire z381_assgn381;
    reg z381_assgn3810;
    reg z186_assgn186;
    wire z7_assgn7;
    wire z9_assgn9;
    wire z11_assgn11;
    wire z395_assgn395;
    reg z395_assgn3950;

    assign x0_0_inp = x0_0;
    assign x1_0_inp = x1_0;
    assign x2_0_inp = x2_0;
    assign x3_0_inp = x3_0;
    assign x0_1_inp = x0_1;
    assign x1_1_inp = x1_1;
    assign x2_1_inp = x2_1;
    assign x3_1_inp = x3_1;
    assign r_inp = r;
    assign L0_0 = (x1_0_inp ^ x2_0_inp);
    assign L1_0 = (x0_0_inp ^ x1_0_inp);
    assign L8_0 = (x2_0_inp ^ x0_0_inp);
    assign L5_0 = (x0_0_inp ^ x3_0_inp);
    assign L0_1 = (x1_1_inp ^ x2_1_inp);
    assign L1_1 = (x0_1_inp ^ x1_1_inp);
    assign L8_1 = (x2_1_inp ^ x0_1_inp);
    assign L5_1 = (x0_1_inp ^ x3_1_inp);
    assign Q0_0 = !L0_0;
    assign Q1_0 = !L1_0;
    assign Q3_0 = !x3_0_inp;
    assign Q4_0 = !x2_0_inp;
    assign Q0_1 = !L0_1;
    assign Q1_1 = !L1_1;
    assign Q3_1 = !x3_1_inp;
    assign Q4_1 = !x2_1_inp;
    assign L2_0 = (Q1_0 ^ x2_0_inp);
    assign L3_0 = (Q0_0 ^ x3_0_inp);
    assign L2_1 = (Q1_1 ^ x2_1_inp);
    assign L3_1 = (Q0_1 ^ x3_1_inp);
    assign p2_domand0 = (Q0_0 & Q1_1);
    assign i1_domand0 = (p2_domand0 ^ r_inp);
    assign p3_domand0 = (Q0_1 & Q1_0);
    assign i2_domand0 = (p3_domand0 ^ r_inp);
    assign p1_domand0 = (Q0_0 & Q1_0);
    assign p4_domand0 = (Q0_1 & Q1_1);
    assign T0_0 = (i1_domand0_reg ^ p1_domand0_reg);
    assign T0_1 = (i2_domand0_reg ^ p4_domand0_reg);
    assign L10_0 = !L2_0;
    assign L10_1 = !L2_1;
    assign p2_domand1 = (x1_0_inp & Q4_1);
    assign i1_domand1 = (p2_domand1 ^ r_inp);
    assign p3_domand1 = (x1_1_inp & Q4_0);
    assign i2_domand1 = (p3_domand1 ^ r_inp);
    assign p1_domand1 = (x1_0_inp & Q4_0);
    assign p4_domand1 = (x1_1_inp & Q4_1);
    assign T2_0 = (i1_domand1_reg ^ p1_domand1_reg);
    assign T2_1 = (i2_domand1_reg ^ p4_domand1_reg);
    assign Q2_0 = (T0_0 ^ L2_0_reg);
    assign L4_0 = (T0_0 ^ T2_0);
    assign Q7_0 = (T0_0 ^ L5_0_reg);
    assign Q6_0 = (L4_0 ^ L3_0_reg);
    assign Q2_1 = (T0_1 ^ L2_1_reg);
    assign L4_1 = (T0_1 ^ T2_1);
    assign Q7_1 = (T0_1 ^ L5_1_reg);
    assign Q6_1 = (L4_1 ^ L3_1_reg);
    assign p2_domand2 = (Q2_0 & Q3_1_reg);
    assign i1_domand2 = (p2_domand2 ^ r_inp_reg);
    assign p3_domand2 = (Q2_1 & Q3_0_reg);
    assign i2_domand2 = (p3_domand2 ^ r_inp_reg);
    assign p1_domand2 = (Q2_0 & Q3_0_reg);
    assign p4_domand2 = (Q2_1 & Q3_1_reg);
    assign T1_0 = (i1_domand2_reg ^ p1_domand2_reg);
    assign T1_1 = (i2_domand2_reg ^ p4_domand2_reg);
    assign p2_domand3 = (Q6_0 & Q7_1);
    assign i1_domand3 = (p2_domand3 ^ r_inp_reg);
    assign p3_domand3 = (Q6_1 & Q7_0);
    assign i2_domand3 = (p3_domand3 ^ r_inp_reg);
    assign p1_domand3 = (Q6_0 & Q7_0);
    assign p4_domand3 = (Q6_1 & Q7_1);
    assign T3_0 = (i1_domand3_reg ^ p1_domand3_reg);
    assign T3_1 = (i2_domand3_reg ^ p4_domand3_reg);
    assign L7_0 = (T0_0_reg ^ T1_0);
    assign z343_assgn343 = L10_0;
    assign L11_0 = (T1_0 ^ z157_assgn157);
    assign L7_1 = (T0_1_reg ^ T1_1);
    assign z349_assgn349 = L10_1;
    assign L11_1 = (T1_1 ^ z161_assgn161);
    assign Y0_01 = (L7_0 ^ T2_0_reg);
    assign z355_assgn355 = L8_0;
    assign Y1_01 = (z166_assgn166 ^ T3_0);
    assign Y0_11 = (L7_1 ^ T2_1_reg);
    assign z361_assgn361 = L8_1;
    assign Y1_11 = (z170_assgn170 ^ T3_1);
    assign z365_assgn365 = x3_0_inp;
    assign z1_assgn1 = (z172_assgn172 ^ Y0_01);
    assign z3_assgn3 = (L11_0 ^ T2_0_reg);
    assign z5_assgn5 = (T2_0 ^ L5_0_reg);
    assign z379_assgn379 = z5_assgn5;
    assign z381_assgn381 = x3_1_inp;
    assign z7_assgn7 = (z186_assgn186 ^ Y0_11);
    assign z9_assgn9 = (L11_1 ^ T2_1_reg);
    assign z11_assgn11 = (T2_1 ^ L5_1_reg);
    assign z395_assgn395 = z11_assgn11;

    always @(posedge clk) begin
        i1_domand0_reg <= i1_domand0;
        p1_domand0_reg <= p1_domand0;
        i2_domand0_reg <= i2_domand0;
        p4_domand0_reg <= p4_domand0;
        i1_domand1_reg <= i1_domand1;
        p1_domand1_reg <= p1_domand1;
        i2_domand1_reg <= i2_domand1;
        p4_domand1_reg <= p4_domand1;
        L2_0_reg <= L2_0;
        L5_0_reg <= L5_0;
        L3_0_reg <= L3_0;
        L2_1_reg <= L2_1;
        L5_1_reg <= L5_1;
        L3_1_reg <= L3_1;
        Q3_1_reg <= Q3_1;
        r_inp_reg <= r_inp;
        Q3_0_reg <= Q3_0;
        i1_domand2_reg <= i1_domand2;
        p1_domand2_reg <= p1_domand2;
        i2_domand2_reg <= i2_domand2;
        p4_domand2_reg <= p4_domand2;
        i1_domand3_reg <= i1_domand3;
        p1_domand3_reg <= p1_domand3;
        i2_domand3_reg <= i2_domand3;
        p4_domand3_reg <= p4_domand3;
        T0_0_reg <= T0_0;
        z343_assgn3430 <= z343_assgn343;
        z157_assgn157 <= z343_assgn3430;
        T0_1_reg <= T0_1;
        z349_assgn3490 <= z349_assgn349;
        z161_assgn161 <= z349_assgn3490;
        T2_0_reg <= T2_0;
        z355_assgn3550 <= z355_assgn355;
        z166_assgn166 <= z355_assgn3550;
        T2_1_reg <= T2_1;
        z361_assgn3610 <= z361_assgn361;
        z170_assgn170 <= z361_assgn3610;
        z365_assgn3650 <= z365_assgn365;
        z172_assgn172 <= z365_assgn3650;
        Y0_0 <= z1_assgn1;
        Y1_0 <= (L7_0 ^ Y1_01);
        Y2_0 <= z3_assgn3;
        z379_assgn3790 <= z379_assgn379;
        Y3_0 <= z379_assgn3790;
        z381_assgn3810 <= z381_assgn381;
        z186_assgn186 <= z381_assgn3810;
        Y0_1 <= z7_assgn7;
        Y1_1 <= (L7_1 ^ Y1_11);
        Y2_1 <= z9_assgn9;
        z395_assgn3950 <= z395_assgn395;
        Y3_1 <= z395_assgn3950;
    end

endmodule

