module sbox(
    clk,
    t0,
    t1,
    r0,
    r1,
    r2,
    r3,
    r4,
    r5,
    dec_0,
    dec_1,
    dec_255,
    dec_169,
    dec_129,
    dec_9,
    dec_72,
    dec_242,
    dec_243,
    dec_152,
    dec_240,
    dec_4,
    dec_15,
    dec_12,
    dec_2,
    dec_3,
    dec_16,
    dec_36,
    dec_220,
    dec_11,
    dec_158,
    dec_45,
    dec_88,
    dec_99,
    y0,
    y1,
);
//INPUTS
    input [7:0] clk;
    input [7:0]  t0;
    input [7:0]  t1;
    input [7:0]  r0;
    input [7:0]  r1;
    input [7:0]  r2;
    input [7:0]  r3;
    input [7:0]  r4;
    input [7:0]  r5;
    input [7:0]  dec_0;
    input [7:0]  dec_1;
    input [7:0]  dec_255;
    input [7:0]  dec_169;
    input [7:0]  dec_129;
    input [7:0]  dec_9;
    input [7:0]  dec_72;
    input [7:0]  dec_242;
    input [7:0]  dec_243;
    input [7:0]  dec_152;
    input [7:0]  dec_240;
    input [7:0]  dec_4;
    input [7:0]  dec_15;
    input [7:0]  dec_12;
    input [7:0]  dec_2;
    input [7:0]  dec_3;
    input [7:0]  dec_16;
    input [7:0]  dec_36;
    input [7:0]  dec_220;
    input [7:0]  dec_11;
    input [7:0]  dec_158;
    input [7:0]  dec_45;
    input [7:0]  dec_88;
    input [7:0]  dec_99;
//OUTPUTS
    output reg [7:0]  y0;
    output reg [7:0]  y1;
//Intermediate values
    wire [7:0] dec_99_inp;
    wire [7:0] dec_88_inp;
    wire [7:0] dec_45_inp;
    wire [7:0] dec_158_inp;
    wire [7:0] dec_11_inp;
    wire [7:0] dec_220_inp;
    wire [7:0] dec_36_inp;
    wire [7:0] dec_16_inp;
    wire [7:0] dec_3_inp;
    wire [7:0] dec_2_inp;
    wire [7:0] dec_12_inp;
    wire [7:0] dec_15_inp;
    wire [7:0] dec_4_inp;
    wire [7:0] dec_240_inp;
    wire [7:0] dec_152_inp;
    wire [7:0] dec_243_inp;
    wire [7:0] dec_242_inp;
    wire [7:0] dec_72_inp;
    wire [7:0] dec_9_inp;
    wire [7:0] dec_129_inp;
    wire [7:0] dec_169_inp;
    wire [7:0] dec_255_inp;
    wire [7:0] dec_1_inp;
    wire [7:0] dec_0_inp;
    wire [7:0] t0_inp;
    wire [7:0] t1_inp;
    wire [7:0] r0_inp;
    wire [7:0] r1_inp;
    wire [7:0] r2_inp;
    wire [7:0] r3_inp;
    wire [7:0] r4_inp;
    wire [7:0] r5_inp;
    wire [7:0] y_G256_newbasis0;
    wire [7:0] tempy1_G256_newbasis0;
    wire [7:0] cond1_G256_newbasis0;
    wire [7:0] negCond1_G256_newbasis0;
    wire [7:0] yxorb1_G256_newbasis0;
    wire [7:0] ny1_G256_newbasis0;
    wire [7:0] tempybooloNegCond1_G256_newbasis0;
    wire [7:0] y1_G256_newbasis0;
    wire [7:0] x1_G256_newbasis0;
    wire [7:0] tempy2_G256_newbasis0;
    wire [7:0] cond2_G256_newbasis0;
    wire [7:0] negCond2_G256_newbasis0;
    wire [7:0] yxorb2_G256_newbasis0;
    wire [7:0] ny2_G256_newbasis0;
    wire [7:0] tempybooloNegCond2_G256_newbasis0;
    wire [7:0] y2_G256_newbasis0;
    wire [7:0] x2_G256_newbasis0;
    wire [7:0] tempy3_G256_newbasis0;
    wire [7:0] cond3_G256_newbasis0;
    wire [7:0] negCond3_G256_newbasis0;
    wire [7:0] yxorb3_G256_newbasis0;
    wire [7:0] ny3_G256_newbasis0;
    wire [7:0] tempybooloNegCond3_G256_newbasis0;
    wire [7:0] y3_G256_newbasis0;
    wire [7:0] x3_G256_newbasis0;
    wire [7:0] tempy4_G256_newbasis0;
    wire [7:0] cond4_G256_newbasis0;
    wire [7:0] negCond4_G256_newbasis0;
    wire [7:0] yxorb4_G256_newbasis0;
    wire [7:0] ny4_G256_newbasis0;
    wire [7:0] tempybooloNegCond4_G256_newbasis0;
    wire [7:0] y4_G256_newbasis0;
    wire [7:0] x4_G256_newbasis0;
    wire [7:0] tempy5_G256_newbasis0;
    wire [7:0] cond5_G256_newbasis0;
    wire [7:0] negCond5_G256_newbasis0;
    wire [7:0] yxorb5_G256_newbasis0;
    wire [7:0] ny5_G256_newbasis0;
    wire [7:0] tempybooloNegCond5_G256_newbasis0;
    wire [7:0] y5_G256_newbasis0;
    wire [7:0] x5_G256_newbasis0;
    wire [7:0] tempy6_G256_newbasis0;
    wire [7:0] cond6_G256_newbasis0;
    wire [7:0] negCond6_G256_newbasis0;
    wire [7:0] yxorb6_G256_newbasis0;
    wire [7:0] ny6_G256_newbasis0;
    wire [7:0] tempybooloNegCond6_G256_newbasis0;
    wire [7:0] y6_G256_newbasis0;
    wire [7:0] x6_G256_newbasis0;
    wire [7:0] tempy7_G256_newbasis0;
    wire [7:0] cond7_G256_newbasis0;
    wire [7:0] negCond7_G256_newbasis0;
    wire [7:0] yxorb7_G256_newbasis0;
    wire [7:0] ny7_G256_newbasis0;
    wire [7:0] tempybooloNegCond7_G256_newbasis0;
    wire [7:0] y7_G256_newbasis0;
    wire [7:0] x7_G256_newbasis0;
    wire [7:0] tempy8_G256_newbasis0;
    wire [7:0] cond8_G256_newbasis0;
    wire [7:0] negCond8_G256_newbasis0;
    wire [7:0] yxorb8_G256_newbasis0;
    wire [7:0] ny8_G256_newbasis0;
    wire [7:0] tempybooloNegCond8_G256_newbasis0;
    wire [7:0] y8_G256_newbasis0;
    wire [7:0] x8_G256_newbasis0;
    wire [7:0] t2;
    wire [7:0] z_y_G256_newbasis0;
    wire [7:0] z_tempy1_G256_newbasis0;
    wire [7:0] z_cond1_G256_newbasis0;
    wire [7:0] z_negCond1_G256_newbasis0;
    wire [7:0] z_yxorb1_G256_newbasis0;
    wire [7:0] z_ny1_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond1_G256_newbasis0;
    wire [7:0] z_y1_G256_newbasis0;
    wire [7:0] z_x1_G256_newbasis0;
    wire [7:0] z_tempy2_G256_newbasis0;
    wire [7:0] z_cond2_G256_newbasis0;
    wire [7:0] z_negCond2_G256_newbasis0;
    wire [7:0] z_yxorb2_G256_newbasis0;
    wire [7:0] z_ny2_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond2_G256_newbasis0;
    wire [7:0] z_y2_G256_newbasis0;
    wire [7:0] z_x2_G256_newbasis0;
    wire [7:0] z_tempy3_G256_newbasis0;
    wire [7:0] z_cond3_G256_newbasis0;
    wire [7:0] z_negCond3_G256_newbasis0;
    wire [7:0] z_yxorb3_G256_newbasis0;
    wire [7:0] z_ny3_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond3_G256_newbasis0;
    wire [7:0] z_y3_G256_newbasis0;
    wire [7:0] z_x3_G256_newbasis0;
    wire [7:0] z_tempy4_G256_newbasis0;
    wire [7:0] z_cond4_G256_newbasis0;
    wire [7:0] z_negCond4_G256_newbasis0;
    wire [7:0] z_yxorb4_G256_newbasis0;
    wire [7:0] z_ny4_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond4_G256_newbasis0;
    wire [7:0] z_y4_G256_newbasis0;
    wire [7:0] z_x4_G256_newbasis0;
    wire [7:0] z_tempy5_G256_newbasis0;
    wire [7:0] z_cond5_G256_newbasis0;
    wire [7:0] z_negCond5_G256_newbasis0;
    wire [7:0] z_yxorb5_G256_newbasis0;
    wire [7:0] z_ny5_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond5_G256_newbasis0;
    wire [7:0] z_y5_G256_newbasis0;
    wire [7:0] z_x5_G256_newbasis0;
    wire [7:0] z_tempy6_G256_newbasis0;
    wire [7:0] z_cond6_G256_newbasis0;
    wire [7:0] z_negCond6_G256_newbasis0;
    wire [7:0] z_yxorb6_G256_newbasis0;
    wire [7:0] z_ny6_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond6_G256_newbasis0;
    wire [7:0] z_y6_G256_newbasis0;
    wire [7:0] z_x6_G256_newbasis0;
    wire [7:0] z_tempy7_G256_newbasis0;
    wire [7:0] z_cond7_G256_newbasis0;
    wire [7:0] z_negCond7_G256_newbasis0;
    wire [7:0] z_yxorb7_G256_newbasis0;
    wire [7:0] z_ny7_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond7_G256_newbasis0;
    wire [7:0] z_y7_G256_newbasis0;
    wire [7:0] z_x7_G256_newbasis0;
    wire [7:0] z_tempy8_G256_newbasis0;
    wire [7:0] z_cond8_G256_newbasis0;
    wire [7:0] z_negCond8_G256_newbasis0;
    wire [7:0] z_yxorb8_G256_newbasis0;
    wire [7:0] z_ny8_G256_newbasis0;
    wire [7:0] z_tempybooloNegCond8_G256_newbasis0;
    wire [7:0] z_y8_G256_newbasis0;
    wire [7:0] z_x8_G256_newbasis0;
    wire [7:0] t3;
    wire [7:0] a0_0_G256_inv0;
    wire [7:0] a1_0_G256_inv0;
    wire [7:0] a0_G256_inv0;
    wire [7:0] a1_G256_inv0;
    wire [7:0] b0_G256_inv0;
    wire [7:0] b1_G256_inv0;
    wire [7:0] a0xorb0_G256_inv0;
    wire [7:0] a1xorb1_G256_inv0;
    wire [7:0] a0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq0_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b0ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] b1ls1_G4_sq1_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_0_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] b1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    wire [7:0] q0_G16_sq_scl0_G256_inv0;
    wire [7:0] q1_G16_sq_scl0_G256_inv0;
    wire [7:0] p0ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] p1ls2_G16_sq_scl0_G256_inv0;
    wire [7:0] c0_G256_inv0;
    wire [7:0] c1_G256_inv0;
    wire [7:0] r00_G16_mul0_G256_inv0;
    wire [7:0] r10_G16_mul0_G256_inv0;
    wire [7:0] r20_G16_mul0_G256_inv0;
    wire [7:0] r30_G16_mul0_G256_inv0;
    wire [7:0] r40_G16_mul0_G256_inv0;
    wire [7:0] r50_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G16_mul0_G256_inv0;
    wire [7:0] a0_G16_mul0_G256_inv0;
    wire [7:0] a1_G16_mul0_G256_inv0;
    wire [7:0] b0_G16_mul0_G256_inv0;
    wire [7:0] b1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G16_mul0_G256_inv0;
    wire [7:0] c0_G16_mul0_G256_inv0;
    wire [7:0] c1_G16_mul0_G256_inv0;
    wire [7:0] d0_G16_mul0_G256_inv0;
    wire [7:0] d1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p1ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul0_G256_inv0;
    wire [7:0] e0_G16_mul0_G256_inv0;
    wire [7:0] e1_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul0_G256_inv0;
    wire [7:0] e01_G16_mul0_G256_inv0;
    wire [7:0] e11_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] e1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p1ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G16_mul0_G256_inv0;
    wire [7:0] p0_G16_mul0_G256_inv0;
    wire [7:0] p1_G16_mul0_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] a1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] b1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] e1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p1ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul0_G256_inv0;
    wire [7:0] q0_0_G16_mul0_G256_inv0;
    wire [7:0] q1_0_G16_mul0_G256_inv0;
    wire [7:0] q0_G16_mul0_G256_inv0;
    wire [7:0] q1_G16_mul0_G256_inv0;
    wire [7:0] p0ls2_G16_mul0_G256_inv0;
    wire [7:0] p1ls2_G16_mul0_G256_inv0;
    wire [7:0] d0_G256_inv0;
    wire [7:0] d1_G256_inv0;
    wire [7:0] c0xord0_G256_inv0;
    wire [7:0] c1xord1_G256_inv0;
    wire [7:0] r00_G16_inv0_G256_inv0;
    wire [7:0] r10_G16_inv0_G256_inv0;
    wire [7:0] r20_G16_inv0_G256_inv0;
    wire [7:0] r30_G16_inv0_G256_inv0;
    wire [7:0] r40_G16_inv0_G256_inv0;
    wire [7:0] r50_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G16_inv0_G256_inv0;
    wire [7:0] a0_G16_inv0_G256_inv0;
    wire [7:0] a1_G16_inv0_G256_inv0;
    wire [7:0] b0_G16_inv0_G256_inv0;
    wire [7:0] b1_G16_inv0_G256_inv0;
    wire [7:0] a0xorb0_G16_inv0_G256_inv0;
    wire [7:0] a1xorb1_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b0ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] b1ls1_G4_sq2_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N1_G16_inv0_G256_inv0;
    wire [7:0] c0_G16_inv0_G256_inv0;
    wire [7:0] c1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] c1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] e1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q1_0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p1ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul3_G16_inv0_G256_inv0;
    wire [7:0] d0_G16_inv0_G256_inv0;
    wire [7:0] d1_G16_inv0_G256_inv0;
    wire [7:0] c0xord0_G16_inv0_G256_inv0;
    wire [7:0] c1xord1_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b0ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] b1ls1_G4_sq3_G16_inv0_G256_inv0;
    wire [7:0] e0_G16_inv0_G256_inv0;
    wire [7:0] e1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] c1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] d1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] e1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q1_0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p1ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul4_G16_inv0_G256_inv0;
    wire [7:0] p0_G16_inv0_G256_inv0;
    wire [7:0] p1_G16_inv0_G256_inv0;
    wire [7:0] r00_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r20_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r30_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r40_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r50_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] a1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] b0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] b1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] c1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] d0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] d1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] axorb_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] cxord_1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m0_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p4_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] e0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] e1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m0_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p4_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r00_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m0_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] m3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p4_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q1_0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p1ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] p0ls1_G4_mul5_G16_inv0_G256_inv0;
    wire [7:0] q0_G16_inv0_G256_inv0;
    wire [7:0] q1_G16_inv0_G256_inv0;
    wire [7:0] p0ls2_G16_inv0_G256_inv0;
    wire [7:0] p1ls2_G16_inv0_G256_inv0;
    wire [7:0] e0_G256_inv0;
    wire [7:0] e1_G256_inv0;
    wire [7:0] r00_G16_mul1_G256_inv0;
    wire [7:0] r10_G16_mul1_G256_inv0;
    wire [7:0] r20_G16_mul1_G256_inv0;
    wire [7:0] r30_G16_mul1_G256_inv0;
    wire [7:0] r40_G16_mul1_G256_inv0;
    wire [7:0] r50_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G16_mul1_G256_inv0;
    wire [7:0] a1_0_G16_mul1_G256_inv0;
    wire [7:0] a0_G16_mul1_G256_inv0;
    wire [7:0] a1_G16_mul1_G256_inv0;
    wire [7:0] b0_G16_mul1_G256_inv0;
    wire [7:0] b1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G16_mul1_G256_inv0;
    wire [7:0] c0_G16_mul1_G256_inv0;
    wire [7:0] c1_G16_mul1_G256_inv0;
    wire [7:0] d0_G16_mul1_G256_inv0;
    wire [7:0] d1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] a1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] b1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m0_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p4_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m0_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p4_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r00_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m0_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] m3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p4_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p1ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul1_G256_inv0;
    wire [7:0] e0_G16_mul1_G256_inv0;
    wire [7:0] e1_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] a1_0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] a1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] b1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul1_G256_inv0;
    wire [7:0] e01_G16_mul1_G256_inv0;
    wire [7:0] e11_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] a1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] b1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m0_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p4_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] e1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m0_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p4_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r00_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m0_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] m3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p4_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p1ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G16_mul1_G256_inv0;
    wire [7:0] p0_G16_mul1_G256_inv0;
    wire [7:0] p1_G16_mul1_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] a1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] b1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m0_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p4_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] e1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m0_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p4_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r00_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m0_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] m3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p4_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p1ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul1_G256_inv0;
    wire [7:0] q0_0_G16_mul1_G256_inv0;
    wire [7:0] q1_0_G16_mul1_G256_inv0;
    wire [7:0] q0_G16_mul1_G256_inv0;
    wire [7:0] q1_G16_mul1_G256_inv0;
    wire [7:0] p0ls2_G16_mul1_G256_inv0;
    wire [7:0] p1ls2_G16_mul1_G256_inv0;
    wire [7:0] p0_G256_inv0;
    wire [7:0] p1_G256_inv0;
    wire [7:0] r00_G16_mul2_G256_inv0;
    wire [7:0] r10_G16_mul2_G256_inv0;
    wire [7:0] r20_G16_mul2_G256_inv0;
    wire [7:0] r30_G16_mul2_G256_inv0;
    wire [7:0] r40_G16_mul2_G256_inv0;
    wire [7:0] r50_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G16_mul2_G256_inv0;
    wire [7:0] a1_0_G16_mul2_G256_inv0;
    wire [7:0] a0_G16_mul2_G256_inv0;
    wire [7:0] a1_G16_mul2_G256_inv0;
    wire [7:0] b0_G16_mul2_G256_inv0;
    wire [7:0] b1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G16_mul2_G256_inv0;
    wire [7:0] c0_G16_mul2_G256_inv0;
    wire [7:0] c1_G16_mul2_G256_inv0;
    wire [7:0] d0_G16_mul2_G256_inv0;
    wire [7:0] d1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] a1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] b1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m0_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p4_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m0_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p4_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r00_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m0_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] m3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p4_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p1ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul0_G16_mul2_G256_inv0;
    wire [7:0] e0_G16_mul2_G256_inv0;
    wire [7:0] e1_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] a1_0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] a1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] b1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p1ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_scl_N0_G16_mul2_G256_inv0;
    wire [7:0] e01_G16_mul2_G256_inv0;
    wire [7:0] e11_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] a1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] b1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m0_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p4_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] e1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m0_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p4_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r00_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m0_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] m3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p4_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p1ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul1_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G16_mul2_G256_inv0;
    wire [7:0] p0_G16_mul2_G256_inv0;
    wire [7:0] p1_G16_mul2_G256_inv0;
    wire [7:0] r00_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r20_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r30_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r40_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r50_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] a1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] b1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] c1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] d1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] axorb_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] cxord_1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m0_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p4_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] e0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] e1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m0_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p4_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r00_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r0_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r1_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r2_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] r3_10_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m0_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] m3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p4_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_1_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_2_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_3_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] y1_4_comar2_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p1ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] p0ls1_G4_mul2_G16_mul2_G256_inv0;
    wire [7:0] q0_0_G16_mul2_G256_inv0;
    wire [7:0] q1_0_G16_mul2_G256_inv0;
    wire [7:0] q0_G16_mul2_G256_inv0;
    wire [7:0] q1_G16_mul2_G256_inv0;
    wire [7:0] p0ls2_G16_mul2_G256_inv0;
    wire [7:0] p1ls2_G16_mul2_G256_inv0;
    wire [7:0] q0_G256_inv0;
    wire [7:0] q1_G256_inv0;
    wire [7:0] p0ls4_G256_inv0;
    wire [7:0] p1ls4_G256_inv0;
    wire [7:0] t4;
    wire [7:0] t5;
    wire [7:0] y_G256_newbasis1;
    wire [7:0] tempy1_G256_newbasis1;
    wire [7:0] cond1_G256_newbasis1;
    wire [7:0] negCond1_G256_newbasis1;
    wire [7:0] yxorb1_G256_newbasis1;
    wire [7:0] ny1_G256_newbasis1;
    wire [7:0] tempybooloNegCond1_G256_newbasis1;
    wire [7:0] y1_G256_newbasis1;
    wire [7:0] x1_G256_newbasis1;
    wire [7:0] tempy2_G256_newbasis1;
    wire [7:0] cond2_G256_newbasis1;
    wire [7:0] negCond2_G256_newbasis1;
    wire [7:0] yxorb2_G256_newbasis1;
    wire [7:0] ny2_G256_newbasis1;
    wire [7:0] tempybooloNegCond2_G256_newbasis1;
    wire [7:0] y2_G256_newbasis1;
    wire [7:0] x2_G256_newbasis1;
    wire [7:0] tempy3_G256_newbasis1;
    wire [7:0] cond3_G256_newbasis1;
    wire [7:0] negCond3_G256_newbasis1;
    wire [7:0] yxorb3_G256_newbasis1;
    wire [7:0] ny3_G256_newbasis1;
    wire [7:0] tempybooloNegCond3_G256_newbasis1;
    wire [7:0] y3_G256_newbasis1;
    wire [7:0] x3_G256_newbasis1;
    wire [7:0] tempy4_G256_newbasis1;
    wire [7:0] cond4_G256_newbasis1;
    wire [7:0] negCond4_G256_newbasis1;
    wire [7:0] yxorb4_G256_newbasis1;
    wire [7:0] ny4_G256_newbasis1;
    wire [7:0] tempybooloNegCond4_G256_newbasis1;
    wire [7:0] y4_G256_newbasis1;
    wire [7:0] x4_G256_newbasis1;
    wire [7:0] tempy5_G256_newbasis1;
    wire [7:0] cond5_G256_newbasis1;
    wire [7:0] negCond5_G256_newbasis1;
    wire [7:0] yxorb5_G256_newbasis1;
    wire [7:0] ny5_G256_newbasis1;
    wire [7:0] tempybooloNegCond5_G256_newbasis1;
    wire [7:0] y5_G256_newbasis1;
    wire [7:0] x5_G256_newbasis1;
    wire [7:0] tempy6_G256_newbasis1;
    wire [7:0] cond6_G256_newbasis1;
    wire [7:0] negCond6_G256_newbasis1;
    wire [7:0] yxorb6_G256_newbasis1;
    wire [7:0] ny6_G256_newbasis1;
    wire [7:0] tempybooloNegCond6_G256_newbasis1;
    wire [7:0] y6_G256_newbasis1;
    wire [7:0] x6_G256_newbasis1;
    wire [7:0] tempy7_G256_newbasis1;
    wire [7:0] cond7_G256_newbasis1;
    wire [7:0] negCond7_G256_newbasis1;
    wire [7:0] yxorb7_G256_newbasis1;
    wire [7:0] ny7_G256_newbasis1;
    wire [7:0] tempybooloNegCond7_G256_newbasis1;
    wire [7:0] y7_G256_newbasis1;
    wire [7:0] x7_G256_newbasis1;
    wire [7:0] tempy8_G256_newbasis1;
    wire [7:0] cond8_G256_newbasis1;
    wire [7:0] negCond8_G256_newbasis1;
    wire [7:0] yxorb8_G256_newbasis1;
    wire [7:0] ny8_G256_newbasis1;
    wire [7:0] tempybooloNegCond8_G256_newbasis1;
    wire [7:0] y8_G256_newbasis1;
    wire [7:0] x8_G256_newbasis1;
    wire [7:0] t6;
    wire [7:0] z_y_G256_newbasis1;
    wire [7:0] z_tempy1_G256_newbasis1;
    wire [7:0] z_cond1_G256_newbasis1;
    wire [7:0] z_negCond1_G256_newbasis1;
    wire [7:0] z_yxorb1_G256_newbasis1;
    wire [7:0] z_ny1_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond1_G256_newbasis1;
    wire [7:0] z_y1_G256_newbasis1;
    wire [7:0] z_x1_G256_newbasis1;
    wire [7:0] z_tempy2_G256_newbasis1;
    wire [7:0] z_cond2_G256_newbasis1;
    wire [7:0] z_negCond2_G256_newbasis1;
    wire [7:0] z_yxorb2_G256_newbasis1;
    wire [7:0] z_ny2_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond2_G256_newbasis1;
    wire [7:0] z_y2_G256_newbasis1;
    wire [7:0] z_x2_G256_newbasis1;
    wire [7:0] z_tempy3_G256_newbasis1;
    wire [7:0] z_cond3_G256_newbasis1;
    wire [7:0] z_negCond3_G256_newbasis1;
    wire [7:0] z_yxorb3_G256_newbasis1;
    wire [7:0] z_ny3_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond3_G256_newbasis1;
    wire [7:0] z_y3_G256_newbasis1;
    wire [7:0] z_x3_G256_newbasis1;
    wire [7:0] z_tempy4_G256_newbasis1;
    wire [7:0] z_cond4_G256_newbasis1;
    wire [7:0] z_negCond4_G256_newbasis1;
    wire [7:0] z_yxorb4_G256_newbasis1;
    wire [7:0] z_ny4_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond4_G256_newbasis1;
    wire [7:0] z_y4_G256_newbasis1;
    wire [7:0] z_x4_G256_newbasis1;
    wire [7:0] z_tempy5_G256_newbasis1;
    wire [7:0] z_cond5_G256_newbasis1;
    wire [7:0] z_negCond5_G256_newbasis1;
    wire [7:0] z_yxorb5_G256_newbasis1;
    wire [7:0] z_ny5_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond5_G256_newbasis1;
    wire [7:0] z_y5_G256_newbasis1;
    wire [7:0] z_x5_G256_newbasis1;
    wire [7:0] z_tempy6_G256_newbasis1;
    wire [7:0] z_cond6_G256_newbasis1;
    wire [7:0] z_negCond6_G256_newbasis1;
    wire [7:0] z_yxorb6_G256_newbasis1;
    wire [7:0] z_ny6_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond6_G256_newbasis1;
    wire [7:0] z_y6_G256_newbasis1;
    wire [7:0] z_x6_G256_newbasis1;
    wire [7:0] z_tempy7_G256_newbasis1;
    wire [7:0] z_cond7_G256_newbasis1;
    wire [7:0] z_negCond7_G256_newbasis1;
    wire [7:0] z_yxorb7_G256_newbasis1;
    wire [7:0] z_ny7_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond7_G256_newbasis1;
    wire [7:0] z_y7_G256_newbasis1;
    wire [7:0] z_x7_G256_newbasis1;
    wire [7:0] z_tempy8_G256_newbasis1;
    wire [7:0] z_cond8_G256_newbasis1;
    wire [7:0] z_negCond8_G256_newbasis1;
    wire [7:0] z_yxorb8_G256_newbasis1;
    wire [7:0] z_ny8_G256_newbasis1;
    wire [7:0] z_tempybooloNegCond8_G256_newbasis1;
    wire [7:0] z_y8_G256_newbasis1;
    wire [7:0] z_x8_G256_newbasis1;
    wire [7:0] t7;

    assign dec_99_inp = dec_99;
    assign dec_88_inp = dec_88;
    assign dec_45_inp = dec_45;
    assign dec_158_inp = dec_158;
    assign dec_11_inp = dec_11;
    assign dec_220_inp = dec_220;
    assign dec_36_inp = dec_36;
    assign dec_16_inp = dec_16;
    assign dec_3_inp = dec_3;
    assign dec_2_inp = dec_2;
    assign dec_12_inp = dec_12;
    assign dec_15_inp = dec_15;
    assign dec_4_inp = dec_4;
    assign dec_240_inp = dec_240;
    assign dec_152_inp = dec_152;
    assign dec_243_inp = dec_243;
    assign dec_242_inp = dec_242;
    assign dec_72_inp = dec_72;
    assign dec_9_inp = dec_9;
    assign dec_129_inp = dec_129;
    assign dec_169_inp = dec_169;
    assign dec_255_inp = dec_255;
    assign dec_1_inp = dec_1;
    assign dec_0_inp = dec_0;
    assign t0_inp = t0;
    assign t1_inp = t1;
    assign r0_inp = r0;
    assign r1_inp = r1;
    assign r2_inp = r2;
    assign r3_inp = r3;
    assign r4_inp = r4;
    assign r5_inp = r5;
    assign y_G256_newbasis0 = dec_0_inp;
    assign tempy1_G256_newbasis0 = y_G256_newbasis0;
    assign cond1_G256_newbasis0 = (t0_inp & dec_1_inp);
    assign negCond1_G256_newbasis0 = !cond1_G256_newbasis0;
    assign yxorb1_G256_newbasis0 = (y_G256_newbasis0 ^ dec_255_inp);
    assign ny1_G256_newbasis0 = (cond1_G256_newbasis0 * yxorb1_G256_newbasis0);
    assign tempybooloNegCond1_G256_newbasis0 = (tempy1_G256_newbasis0 * negCond1_G256_newbasis0);
    assign y1_G256_newbasis0 = (ny1_G256_newbasis0 + tempybooloNegCond1_G256_newbasis0);
    assign x1_G256_newbasis0 = (t0_inp >> dec_1_inp);
    assign tempy2_G256_newbasis0 = y1_G256_newbasis0;
    assign cond2_G256_newbasis0 = (x1_G256_newbasis0 & dec_1_inp);
    assign negCond2_G256_newbasis0 = !cond2_G256_newbasis0;
    assign yxorb2_G256_newbasis0 = (y1_G256_newbasis0 ^ dec_169_inp);
    assign ny2_G256_newbasis0 = (cond2_G256_newbasis0 * yxorb2_G256_newbasis0);
    assign tempybooloNegCond2_G256_newbasis0 = (tempy2_G256_newbasis0 * negCond2_G256_newbasis0);
    assign y2_G256_newbasis0 = (ny2_G256_newbasis0 + tempybooloNegCond2_G256_newbasis0);
    assign x2_G256_newbasis0 = (x1_G256_newbasis0 >> dec_1_inp);
    assign tempy3_G256_newbasis0 = y2_G256_newbasis0;
    assign cond3_G256_newbasis0 = (x2_G256_newbasis0 & dec_1_inp);
    assign negCond3_G256_newbasis0 = !cond3_G256_newbasis0;
    assign yxorb3_G256_newbasis0 = (y2_G256_newbasis0 ^ dec_129_inp);
    assign ny3_G256_newbasis0 = (cond3_G256_newbasis0 * yxorb3_G256_newbasis0);
    assign tempybooloNegCond3_G256_newbasis0 = (tempy3_G256_newbasis0 * negCond3_G256_newbasis0);
    assign y3_G256_newbasis0 = (ny3_G256_newbasis0 + tempybooloNegCond3_G256_newbasis0);
    assign x3_G256_newbasis0 = (x2_G256_newbasis0 >> dec_1_inp);
    assign tempy4_G256_newbasis0 = y3_G256_newbasis0;
    assign cond4_G256_newbasis0 = (x3_G256_newbasis0 & dec_1_inp);
    assign negCond4_G256_newbasis0 = !cond4_G256_newbasis0;
    assign yxorb4_G256_newbasis0 = (y3_G256_newbasis0 ^ dec_9_inp);
    assign ny4_G256_newbasis0 = (cond4_G256_newbasis0 * yxorb4_G256_newbasis0);
    assign tempybooloNegCond4_G256_newbasis0 = (tempy4_G256_newbasis0 * negCond4_G256_newbasis0);
    assign y4_G256_newbasis0 = (ny4_G256_newbasis0 + tempybooloNegCond4_G256_newbasis0);
    assign x4_G256_newbasis0 = (x3_G256_newbasis0 >> dec_1_inp);
    assign tempy5_G256_newbasis0 = y4_G256_newbasis0;
    assign cond5_G256_newbasis0 = (x4_G256_newbasis0 & dec_1_inp);
    assign negCond5_G256_newbasis0 = !cond5_G256_newbasis0;
    assign yxorb5_G256_newbasis0 = (y4_G256_newbasis0 ^ dec_72_inp);
    assign ny5_G256_newbasis0 = (cond5_G256_newbasis0 * yxorb5_G256_newbasis0);
    assign tempybooloNegCond5_G256_newbasis0 = (tempy5_G256_newbasis0 * negCond5_G256_newbasis0);
    assign y5_G256_newbasis0 = (ny5_G256_newbasis0 + tempybooloNegCond5_G256_newbasis0);
    assign x5_G256_newbasis0 = (x4_G256_newbasis0 >> dec_1_inp);
    assign tempy6_G256_newbasis0 = y5_G256_newbasis0;
    assign cond6_G256_newbasis0 = (x5_G256_newbasis0 & dec_1_inp);
    assign negCond6_G256_newbasis0 = !cond6_G256_newbasis0;
    assign yxorb6_G256_newbasis0 = (y5_G256_newbasis0 ^ dec_242_inp);
    assign ny6_G256_newbasis0 = (cond6_G256_newbasis0 * yxorb6_G256_newbasis0);
    assign tempybooloNegCond6_G256_newbasis0 = (tempy6_G256_newbasis0 * negCond6_G256_newbasis0);
    assign y6_G256_newbasis0 = (ny6_G256_newbasis0 + tempybooloNegCond6_G256_newbasis0);
    assign x6_G256_newbasis0 = (x5_G256_newbasis0 >> dec_1_inp);
    assign tempy7_G256_newbasis0 = y6_G256_newbasis0;
    assign cond7_G256_newbasis0 = (x6_G256_newbasis0 & dec_1_inp);
    assign negCond7_G256_newbasis0 = !cond7_G256_newbasis0;
    assign yxorb7_G256_newbasis0 = (y6_G256_newbasis0 ^ dec_243_inp);
    assign ny7_G256_newbasis0 = (cond7_G256_newbasis0 * yxorb7_G256_newbasis0);
    assign tempybooloNegCond7_G256_newbasis0 = (tempy7_G256_newbasis0 * negCond7_G256_newbasis0);
    assign y7_G256_newbasis0 = (ny7_G256_newbasis0 + tempybooloNegCond7_G256_newbasis0);
    assign x7_G256_newbasis0 = (x6_G256_newbasis0 >> dec_1_inp);
    assign tempy8_G256_newbasis0 = y7_G256_newbasis0;
    assign cond8_G256_newbasis0 = (x7_G256_newbasis0 & dec_1_inp);
    assign negCond8_G256_newbasis0 = !cond8_G256_newbasis0;
    assign yxorb8_G256_newbasis0 = (y7_G256_newbasis0 ^ dec_152_inp);
    assign ny8_G256_newbasis0 = (cond8_G256_newbasis0 * yxorb8_G256_newbasis0);
    assign tempybooloNegCond8_G256_newbasis0 = (tempy8_G256_newbasis0 * negCond8_G256_newbasis0);
    assign y8_G256_newbasis0 = (ny8_G256_newbasis0 + tempybooloNegCond8_G256_newbasis0);
    assign x8_G256_newbasis0 = (x7_G256_newbasis0 >> dec_1_inp);
    assign t2 = y8_G256_newbasis0;
    assign z_y_G256_newbasis0 = dec_0_inp;
    assign z_tempy1_G256_newbasis0 = z_y_G256_newbasis0;
    assign z_cond1_G256_newbasis0 = (t1_inp & dec_1_inp);
    assign z_negCond1_G256_newbasis0 = !z_cond1_G256_newbasis0;
    assign z_yxorb1_G256_newbasis0 = (z_y_G256_newbasis0 ^ dec_255_inp);
    assign z_ny1_G256_newbasis0 = (z_cond1_G256_newbasis0 * z_yxorb1_G256_newbasis0);
    assign z_tempybooloNegCond1_G256_newbasis0 = (z_tempy1_G256_newbasis0 * z_negCond1_G256_newbasis0);
    assign z_y1_G256_newbasis0 = (z_ny1_G256_newbasis0 + z_tempybooloNegCond1_G256_newbasis0);
    assign z_x1_G256_newbasis0 = (t1_inp >> dec_1_inp);
    assign z_tempy2_G256_newbasis0 = z_y1_G256_newbasis0;
    assign z_cond2_G256_newbasis0 = (z_x1_G256_newbasis0 & dec_1_inp);
    assign z_negCond2_G256_newbasis0 = !z_cond2_G256_newbasis0;
    assign z_yxorb2_G256_newbasis0 = (z_y1_G256_newbasis0 ^ dec_169_inp);
    assign z_ny2_G256_newbasis0 = (z_cond2_G256_newbasis0 * z_yxorb2_G256_newbasis0);
    assign z_tempybooloNegCond2_G256_newbasis0 = (z_tempy2_G256_newbasis0 * z_negCond2_G256_newbasis0);
    assign z_y2_G256_newbasis0 = (z_ny2_G256_newbasis0 + z_tempybooloNegCond2_G256_newbasis0);
    assign z_x2_G256_newbasis0 = (z_x1_G256_newbasis0 >> dec_1_inp);
    assign z_tempy3_G256_newbasis0 = z_y2_G256_newbasis0;
    assign z_cond3_G256_newbasis0 = (z_x2_G256_newbasis0 & dec_1_inp);
    assign z_negCond3_G256_newbasis0 = !z_cond3_G256_newbasis0;
    assign z_yxorb3_G256_newbasis0 = (z_y2_G256_newbasis0 ^ dec_129_inp);
    assign z_ny3_G256_newbasis0 = (z_cond3_G256_newbasis0 * z_yxorb3_G256_newbasis0);
    assign z_tempybooloNegCond3_G256_newbasis0 = (z_tempy3_G256_newbasis0 * z_negCond3_G256_newbasis0);
    assign z_y3_G256_newbasis0 = (z_ny3_G256_newbasis0 + z_tempybooloNegCond3_G256_newbasis0);
    assign z_x3_G256_newbasis0 = (z_x2_G256_newbasis0 >> dec_1_inp);
    assign z_tempy4_G256_newbasis0 = z_y3_G256_newbasis0;
    assign z_cond4_G256_newbasis0 = (z_x3_G256_newbasis0 & dec_1_inp);
    assign z_negCond4_G256_newbasis0 = !z_cond4_G256_newbasis0;
    assign z_yxorb4_G256_newbasis0 = (z_y3_G256_newbasis0 ^ dec_9_inp);
    assign z_ny4_G256_newbasis0 = (z_cond4_G256_newbasis0 * z_yxorb4_G256_newbasis0);
    assign z_tempybooloNegCond4_G256_newbasis0 = (z_tempy4_G256_newbasis0 * z_negCond4_G256_newbasis0);
    assign z_y4_G256_newbasis0 = (z_ny4_G256_newbasis0 + z_tempybooloNegCond4_G256_newbasis0);
    assign z_x4_G256_newbasis0 = (z_x3_G256_newbasis0 >> dec_1_inp);
    assign z_tempy5_G256_newbasis0 = z_y4_G256_newbasis0;
    assign z_cond5_G256_newbasis0 = (z_x4_G256_newbasis0 & dec_1_inp);
    assign z_negCond5_G256_newbasis0 = !z_cond5_G256_newbasis0;
    assign z_yxorb5_G256_newbasis0 = (z_y4_G256_newbasis0 ^ dec_72_inp);
    assign z_ny5_G256_newbasis0 = (z_cond5_G256_newbasis0 * z_yxorb5_G256_newbasis0);
    assign z_tempybooloNegCond5_G256_newbasis0 = (z_tempy5_G256_newbasis0 * z_negCond5_G256_newbasis0);
    assign z_y5_G256_newbasis0 = (z_ny5_G256_newbasis0 + z_tempybooloNegCond5_G256_newbasis0);
    assign z_x5_G256_newbasis0 = (z_x4_G256_newbasis0 >> dec_1_inp);
    assign z_tempy6_G256_newbasis0 = z_y5_G256_newbasis0;
    assign z_cond6_G256_newbasis0 = (z_x5_G256_newbasis0 & dec_1_inp);
    assign z_negCond6_G256_newbasis0 = !z_cond6_G256_newbasis0;
    assign z_yxorb6_G256_newbasis0 = (z_y5_G256_newbasis0 ^ dec_242_inp);
    assign z_ny6_G256_newbasis0 = (z_cond6_G256_newbasis0 * z_yxorb6_G256_newbasis0);
    assign z_tempybooloNegCond6_G256_newbasis0 = (z_tempy6_G256_newbasis0 * z_negCond6_G256_newbasis0);
    assign z_y6_G256_newbasis0 = (z_ny6_G256_newbasis0 + z_tempybooloNegCond6_G256_newbasis0);
    assign z_x6_G256_newbasis0 = (z_x5_G256_newbasis0 >> dec_1_inp);
    assign z_tempy7_G256_newbasis0 = z_y6_G256_newbasis0;
    assign z_cond7_G256_newbasis0 = (z_x6_G256_newbasis0 & dec_1_inp);
    assign z_negCond7_G256_newbasis0 = !z_cond7_G256_newbasis0;
    assign z_yxorb7_G256_newbasis0 = (z_y6_G256_newbasis0 ^ dec_243_inp);
    assign z_ny7_G256_newbasis0 = (z_cond7_G256_newbasis0 * z_yxorb7_G256_newbasis0);
    assign z_tempybooloNegCond7_G256_newbasis0 = (z_tempy7_G256_newbasis0 * z_negCond7_G256_newbasis0);
    assign z_y7_G256_newbasis0 = (z_ny7_G256_newbasis0 + z_tempybooloNegCond7_G256_newbasis0);
    assign z_x7_G256_newbasis0 = (z_x6_G256_newbasis0 >> dec_1_inp);
    assign z_tempy8_G256_newbasis0 = z_y7_G256_newbasis0;
    assign z_cond8_G256_newbasis0 = (z_x7_G256_newbasis0 & dec_1_inp);
    assign z_negCond8_G256_newbasis0 = !z_cond8_G256_newbasis0;
    assign z_yxorb8_G256_newbasis0 = (z_y7_G256_newbasis0 ^ dec_152_inp);
    assign z_ny8_G256_newbasis0 = (z_cond8_G256_newbasis0 * z_yxorb8_G256_newbasis0);
    assign z_tempybooloNegCond8_G256_newbasis0 = (z_tempy8_G256_newbasis0 * z_negCond8_G256_newbasis0);
    assign z_y8_G256_newbasis0 = (z_ny8_G256_newbasis0 + z_tempybooloNegCond8_G256_newbasis0);
    assign z_x8_G256_newbasis0 = (z_x7_G256_newbasis0 >> dec_1_inp);
    assign t3 = z_y8_G256_newbasis0;
    assign a0_0_G256_inv0 = (t2 & dec_240_inp);
    assign a1_0_G256_inv0 = (t3 & dec_240_inp);
    assign a0_G256_inv0 = (a0_0_G256_inv0 >> dec_4_inp);
    assign a1_G256_inv0 = (a1_0_G256_inv0 >> dec_4_inp);
    assign b0_G256_inv0 = (t2 & dec_15_inp);
    assign b1_G256_inv0 = (t3 & dec_15_inp);
    assign a0xorb0_G256_inv0 = (a0_G256_inv0 ^ b0_G256_inv0);
    assign a1xorb1_G256_inv0 = (a1_G256_inv0 ^ b1_G256_inv0);
    assign a0_0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_12_inp);
    assign a0_G16_sq_scl0_G256_inv0 = (a0_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign a1_G16_sq_scl0_G256_inv0 = (a1_0_G16_sq_scl0_G256_inv0 >> dec_2_inp);
    assign b0_G16_sq_scl0_G256_inv0 = (a0xorb0_G256_inv0 & dec_3_inp);
    assign b1_G16_sq_scl0_G256_inv0 = (a1xorb1_G256_inv0 & dec_3_inp);
    assign p0_0_G16_sq_scl0_G256_inv0 = (a0_G16_sq_scl0_G256_inv0 ^ b0_G16_sq_scl0_G256_inv0);
    assign p1_0_G16_sq_scl0_G256_inv0 = (a1_G16_sq_scl0_G256_inv0 ^ b1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq0_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq0_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq0_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq0_G16_sq_scl0_G256_inv0 = (p0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq0_G16_sq_scl0_G256_inv0 = (p1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b0_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 = (b1_G4_sq0_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a0_G4_sq0_G16_sq_scl0_G256_inv0);
    assign p1_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq0_G16_sq_scl0_G256_inv0 | a1_G4_sq0_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq1_G16_sq_scl0_G256_inv0 = (a0_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq1_G16_sq_scl0_G256_inv0 = (a1_0_G4_sq1_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b0_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 = (b1_G4_sq1_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_sq_scl0_G256_inv0 = (b0ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a0_G4_sq1_G16_sq_scl0_G256_inv0);
    assign q1_0_G16_sq_scl0_G256_inv0 = (b1ls1_G4_sq1_G16_sq_scl0_G256_inv0 | a1_G4_sq1_G16_sq_scl0_G256_inv0);
    assign a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_0_G4_scl_N20_G16_sq_scl0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q0_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (q1_0_G16_sq_scl0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a0_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (a1_G4_scl_N20_G16_sq_scl0_G256_inv0 ^ b1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q0_G4_scl_N20_G16_sq_scl0_G256_inv0 = a0_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign q1_G4_scl_N20_G16_sq_scl0_G256_inv0 = a1_G4_scl_N20_G16_sq_scl0_G256_inv0;
    assign p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p1_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 = (p0_G4_scl_N20_G16_sq_scl0_G256_inv0 << dec_1_inp);
    assign q0_G16_sq_scl0_G256_inv0 = (p0ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q0_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign q1_G16_sq_scl0_G256_inv0 = (p1ls1_G4_scl_N20_G16_sq_scl0_G256_inv0 | q1_G4_scl_N20_G16_sq_scl0_G256_inv0);
    assign p0ls2_G16_sq_scl0_G256_inv0 = (p0_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_sq_scl0_G256_inv0 = (p1_G16_sq_scl0_G256_inv0 << dec_2_inp);
    assign c0_G256_inv0 = (p0ls2_G16_sq_scl0_G256_inv0 | q0_G16_sq_scl0_G256_inv0);
    assign c1_G256_inv0 = (p1ls2_G16_sq_scl0_G256_inv0 | q1_G16_sq_scl0_G256_inv0);
    assign r00_G16_mul0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul0_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul0_G256_inv0 = (a0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul0_G256_inv0 = (a1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul0_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul0_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul0_G256_inv0 = (c0_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul0_G256_inv0 = (c1_0_G16_mul0_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul0_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul0_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 ^ b0_G16_mul0_G256_inv0);
    assign cxord_0_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 ^ d0_G16_mul0_G256_inv0);
    assign axorb_1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 ^ b1_G16_mul0_G256_inv0);
    assign cxord_1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 ^ d1_G16_mul0_G256_inv0);
    assign r00_G4_mul0_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul0_G256_inv0 = (a0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul0_G256_inv0 = (a1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul0_G256_inv0 = (c0_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul0_G256_inv0 = (c1_0_G4_mul0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ b0_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ d0_G4_mul0_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ b1_G4_mul0_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ d1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul0_G256_inv0 = (axorb_0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul0_G256_inv0 = (cxord_1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul0_G256_inv0 = (cxord_0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul0_G16_mul0_G256_inv0 = (axorb_1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul0_G16_mul0_G256_inv0 = (m0_comar0_G4_mul0_G16_mul0_G256_inv0 & m1_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign p3_comar0_G4_mul0_G16_mul0_G256_inv0 = (m3_comar0_G4_mul0_G16_mul0_G256_inv0 & m2_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_comar0_G4_mul0_G16_mul0_G256_inv0 = (m0_comar0_G4_mul0_G16_mul0_G256_inv0 & m2_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign p4_comar0_G4_mul0_G16_mul0_G256_inv0 = (m3_comar0_G4_mul0_G16_mul0_G256_inv0 & m1_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i0_comar0_G4_mul0_G16_mul0_G256_inv0 = (p1_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i1_comar0_G4_mul0_G16_mul0_G256_inv0 = (p2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i2_comar0_G4_mul0_G16_mul0_G256_inv0 = (p3_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i3_comar0_G4_mul0_G16_mul0_G256_inv0 = (p4_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0 = (i1_comar0_G4_mul0_G16_mul0_G256_inv0 ^ i2_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0 = (i0_comar0_G4_mul0_G16_mul0_G256_inv0 ^ i3_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign e0_G4_mul0_G16_mul0_G256_inv0 = (i1xori2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_1_comar0_G4_mul0_G16_mul0_G256_inv0 = (r00_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul0_G256_inv0 = (a0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul0_G256_inv0 = (c1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul0_G256_inv0 = (c0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul0_G16_mul0_G256_inv0 = (a1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul0_G16_mul0_G256_inv0 = (m0_comar1_G4_mul0_G16_mul0_G256_inv0 & m1_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p3_comar1_G4_mul0_G16_mul0_G256_inv0 = (m3_comar1_G4_mul0_G16_mul0_G256_inv0 & m2_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p1_comar1_G4_mul0_G16_mul0_G256_inv0 = (m0_comar1_G4_mul0_G16_mul0_G256_inv0 & m2_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p4_comar1_G4_mul0_G16_mul0_G256_inv0 = (m3_comar1_G4_mul0_G16_mul0_G256_inv0 & m1_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i0_comar1_G4_mul0_G16_mul0_G256_inv0 = (p1_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i1_comar1_G4_mul0_G16_mul0_G256_inv0 = (p2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i2_comar1_G4_mul0_G16_mul0_G256_inv0 = (p3_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i3_comar1_G4_mul0_G16_mul0_G256_inv0 = (p4_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0 = (i1_comar1_G4_mul0_G16_mul0_G256_inv0 ^ i2_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0 = (i0_comar1_G4_mul0_G16_mul0_G256_inv0 ^ i3_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p0_0_G4_mul0_G16_mul0_G256_inv0 = (i1xori2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_1_comar1_G4_mul0_G16_mul0_G256_inv0 = (r00_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p1_0_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul0_G256_inv0);
    assign p0_G4_mul0_G16_mul0_G256_inv0 = (p0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign p1_G4_mul0_G16_mul0_G256_inv0 = (p1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul0_G256_inv0 = (r00_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r10_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r20_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r30_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r40_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul0_G256_inv0 = (r50_G4_mul0_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul0_G256_inv0 = (b0_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul0_G256_inv0 = (d1_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul0_G256_inv0 = (d0_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul0_G16_mul0_G256_inv0 = (b1_G4_mul0_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul0_G16_mul0_G256_inv0 = (m0_comar2_G4_mul0_G16_mul0_G256_inv0 & m1_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign p3_comar2_G4_mul0_G16_mul0_G256_inv0 = (m3_comar2_G4_mul0_G16_mul0_G256_inv0 & m2_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign p1_comar2_G4_mul0_G16_mul0_G256_inv0 = (m0_comar2_G4_mul0_G16_mul0_G256_inv0 & m2_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign p4_comar2_G4_mul0_G16_mul0_G256_inv0 = (m3_comar2_G4_mul0_G16_mul0_G256_inv0 & m1_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i0_comar2_G4_mul0_G16_mul0_G256_inv0 = (p1_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i1_comar2_G4_mul0_G16_mul0_G256_inv0 = (p2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i2_comar2_G4_mul0_G16_mul0_G256_inv0 = (p3_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i3_comar2_G4_mul0_G16_mul0_G256_inv0 = (p4_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0 = (i1_comar2_G4_mul0_G16_mul0_G256_inv0 ^ i2_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0 = (i0_comar2_G4_mul0_G16_mul0_G256_inv0 ^ i3_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign q0_0_G4_mul0_G16_mul0_G256_inv0 = (i1xori2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_1_comar2_G4_mul0_G16_mul0_G256_inv0 = (r00_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign q1_0_G4_mul0_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul0_G256_inv0);
    assign q0_G4_mul0_G16_mul0_G256_inv0 = (q0_0_G4_mul0_G16_mul0_G256_inv0 ^ e0_G4_mul0_G16_mul0_G256_inv0);
    assign q1_G4_mul0_G16_mul0_G256_inv0 = (q1_0_G4_mul0_G16_mul0_G256_inv0 ^ e1_G4_mul0_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul0_G256_inv0 = (p1_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul0_G16_mul0_G256_inv0 = (p0_G4_mul0_G16_mul0_G256_inv0 << dec_1_inp);
    assign e0_G16_mul0_G256_inv0 = (p1ls1_G4_mul0_G16_mul0_G256_inv0 | q1_G4_mul0_G16_mul0_G256_inv0);
    assign e1_G16_mul0_G256_inv0 = (p0ls1_G4_mul0_G16_mul0_G256_inv0 | q0_G4_mul0_G16_mul0_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_0_G4_scl_N0_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul0_G256_inv0 = (e0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N0_G16_mul0_G256_inv0 = (e1_G16_mul0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul0_G256_inv0 = b0_G4_scl_N0_G16_mul0_G256_inv0;
    assign p1_G4_scl_N0_G16_mul0_G256_inv0 = b1_G4_scl_N0_G16_mul0_G256_inv0;
    assign q0_G4_scl_N0_G16_mul0_G256_inv0 = (a0_G4_scl_N0_G16_mul0_G256_inv0 ^ b0_G4_scl_N0_G16_mul0_G256_inv0);
    assign q1_G4_scl_N0_G16_mul0_G256_inv0 = (a1_G4_scl_N0_G16_mul0_G256_inv0 ^ b1_G4_scl_N0_G16_mul0_G256_inv0);
    assign p1ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p1_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N0_G16_mul0_G256_inv0 = (p0_G4_scl_N0_G16_mul0_G256_inv0 << dec_1_inp);
    assign e01_G16_mul0_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul0_G256_inv0 | q0_G4_scl_N0_G16_mul0_G256_inv0);
    assign e11_G16_mul0_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul0_G256_inv0 | q1_G4_scl_N0_G16_mul0_G256_inv0);
    assign r00_G4_mul1_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul0_G256_inv0 = (a0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul0_G256_inv0 = (a1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul0_G256_inv0 = (a0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul0_G256_inv0 = (a1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul0_G256_inv0 = (c0_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul0_G256_inv0 = (c1_0_G4_mul1_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul0_G256_inv0 = (c0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul0_G256_inv0 = (c1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ b0_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ d0_G4_mul1_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ b1_G4_mul1_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ d1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul0_G256_inv0 = (axorb_0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul0_G256_inv0 = (cxord_1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul0_G256_inv0 = (cxord_0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul1_G16_mul0_G256_inv0 = (axorb_1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul1_G16_mul0_G256_inv0 = (m0_comar0_G4_mul1_G16_mul0_G256_inv0 & m1_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign p3_comar0_G4_mul1_G16_mul0_G256_inv0 = (m3_comar0_G4_mul1_G16_mul0_G256_inv0 & m2_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_comar0_G4_mul1_G16_mul0_G256_inv0 = (m0_comar0_G4_mul1_G16_mul0_G256_inv0 & m2_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign p4_comar0_G4_mul1_G16_mul0_G256_inv0 = (m3_comar0_G4_mul1_G16_mul0_G256_inv0 & m1_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i0_comar0_G4_mul1_G16_mul0_G256_inv0 = (p1_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i1_comar0_G4_mul1_G16_mul0_G256_inv0 = (p2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i2_comar0_G4_mul1_G16_mul0_G256_inv0 = (p3_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i3_comar0_G4_mul1_G16_mul0_G256_inv0 = (p4_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0 = (i1_comar0_G4_mul1_G16_mul0_G256_inv0 ^ i2_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0 = (i0_comar0_G4_mul1_G16_mul0_G256_inv0 ^ i3_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign e0_G4_mul1_G16_mul0_G256_inv0 = (i1xori2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_1_comar0_G4_mul1_G16_mul0_G256_inv0 = (r00_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign e1_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul0_G256_inv0 = (a0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul0_G256_inv0 = (c1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul0_G256_inv0 = (c0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul1_G16_mul0_G256_inv0 = (a1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul1_G16_mul0_G256_inv0 = (m0_comar1_G4_mul1_G16_mul0_G256_inv0 & m1_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p3_comar1_G4_mul1_G16_mul0_G256_inv0 = (m3_comar1_G4_mul1_G16_mul0_G256_inv0 & m2_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_comar1_G4_mul1_G16_mul0_G256_inv0 = (m0_comar1_G4_mul1_G16_mul0_G256_inv0 & m2_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p4_comar1_G4_mul1_G16_mul0_G256_inv0 = (m3_comar1_G4_mul1_G16_mul0_G256_inv0 & m1_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i0_comar1_G4_mul1_G16_mul0_G256_inv0 = (p1_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i1_comar1_G4_mul1_G16_mul0_G256_inv0 = (p2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i2_comar1_G4_mul1_G16_mul0_G256_inv0 = (p3_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i3_comar1_G4_mul1_G16_mul0_G256_inv0 = (p4_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0 = (i1_comar1_G4_mul1_G16_mul0_G256_inv0 ^ i2_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0 = (i0_comar1_G4_mul1_G16_mul0_G256_inv0 ^ i3_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p0_0_G4_mul1_G16_mul0_G256_inv0 = (i1xori2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_1_comar1_G4_mul1_G16_mul0_G256_inv0 = (r00_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G4_mul1_G16_mul0_G256_inv0 = (p0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign p1_G4_mul1_G16_mul0_G256_inv0 = (p1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul0_G256_inv0 = (r00_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r10_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r20_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r30_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r40_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul0_G256_inv0 = (r50_G4_mul1_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul0_G256_inv0 = (b0_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul0_G256_inv0 = (d1_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul0_G256_inv0 = (d0_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul1_G16_mul0_G256_inv0 = (b1_G4_mul1_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul1_G16_mul0_G256_inv0 = (m0_comar2_G4_mul1_G16_mul0_G256_inv0 & m1_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign p3_comar2_G4_mul1_G16_mul0_G256_inv0 = (m3_comar2_G4_mul1_G16_mul0_G256_inv0 & m2_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign p1_comar2_G4_mul1_G16_mul0_G256_inv0 = (m0_comar2_G4_mul1_G16_mul0_G256_inv0 & m2_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign p4_comar2_G4_mul1_G16_mul0_G256_inv0 = (m3_comar2_G4_mul1_G16_mul0_G256_inv0 & m1_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i0_comar2_G4_mul1_G16_mul0_G256_inv0 = (p1_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i1_comar2_G4_mul1_G16_mul0_G256_inv0 = (p2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i2_comar2_G4_mul1_G16_mul0_G256_inv0 = (p3_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i3_comar2_G4_mul1_G16_mul0_G256_inv0 = (p4_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0 = (i1_comar2_G4_mul1_G16_mul0_G256_inv0 ^ i2_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0 = (i0_comar2_G4_mul1_G16_mul0_G256_inv0 ^ i3_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign q0_0_G4_mul1_G16_mul0_G256_inv0 = (i1xori2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_1_comar2_G4_mul1_G16_mul0_G256_inv0 = (r00_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign q1_0_G4_mul1_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul0_G256_inv0);
    assign q0_G4_mul1_G16_mul0_G256_inv0 = (q0_0_G4_mul1_G16_mul0_G256_inv0 ^ e0_G4_mul1_G16_mul0_G256_inv0);
    assign q1_G4_mul1_G16_mul0_G256_inv0 = (q1_0_G4_mul1_G16_mul0_G256_inv0 ^ e1_G4_mul1_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul0_G256_inv0 = (p1_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul1_G16_mul0_G256_inv0 = (p0_G4_mul1_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul1_G16_mul0_G256_inv0 | q1_G4_mul1_G16_mul0_G256_inv0);
    assign p1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul1_G16_mul0_G256_inv0 | q0_G4_mul1_G16_mul0_G256_inv0);
    assign p0_G16_mul0_G256_inv0 = (p0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign p1_G16_mul0_G256_inv0 = (p1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign r00_G4_mul2_G16_mul0_G256_inv0 = (r00_G16_mul0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul0_G256_inv0 = (r10_G16_mul0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul0_G256_inv0 = (r20_G16_mul0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul0_G256_inv0 = (r30_G16_mul0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul0_G256_inv0 = (r40_G16_mul0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul0_G256_inv0 = (r50_G16_mul0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul0_G256_inv0 = (a0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul0_G256_inv0 = (a1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul0_G256_inv0 = (b0_G16_mul0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul0_G256_inv0 = (b1_G16_mul0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul0_G256_inv0 = (c0_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul0_G256_inv0 = (c1_0_G4_mul2_G16_mul0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul0_G256_inv0 = (d0_G16_mul0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul0_G256_inv0 = (d1_G16_mul0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ b0_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ d0_G4_mul2_G16_mul0_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ b1_G4_mul2_G16_mul0_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ d1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul0_G256_inv0 = (axorb_0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul0_G256_inv0 = (cxord_1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul0_G256_inv0 = (cxord_0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar0_G4_mul2_G16_mul0_G256_inv0 = (axorb_1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar0_G4_mul2_G16_mul0_G256_inv0 = (m0_comar0_G4_mul2_G16_mul0_G256_inv0 & m1_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign p3_comar0_G4_mul2_G16_mul0_G256_inv0 = (m3_comar0_G4_mul2_G16_mul0_G256_inv0 & m2_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_comar0_G4_mul2_G16_mul0_G256_inv0 = (m0_comar0_G4_mul2_G16_mul0_G256_inv0 & m2_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign p4_comar0_G4_mul2_G16_mul0_G256_inv0 = (m3_comar0_G4_mul2_G16_mul0_G256_inv0 & m1_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i0_comar0_G4_mul2_G16_mul0_G256_inv0 = (p1_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i1_comar0_G4_mul2_G16_mul0_G256_inv0 = (p2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i2_comar0_G4_mul2_G16_mul0_G256_inv0 = (p3_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i3_comar0_G4_mul2_G16_mul0_G256_inv0 = (p4_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0 = (i1_comar0_G4_mul2_G16_mul0_G256_inv0 ^ i2_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0 = (i0_comar0_G4_mul2_G16_mul0_G256_inv0 ^ i3_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign e0_G4_mul2_G16_mul0_G256_inv0 = (i1xori2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_1_comar0_G4_mul2_G16_mul0_G256_inv0 = (r00_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign e1_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul0_G256_inv0 = (a0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul0_G256_inv0 = (c1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul0_G256_inv0 = (c0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar1_G4_mul2_G16_mul0_G256_inv0 = (a1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar1_G4_mul2_G16_mul0_G256_inv0 = (m0_comar1_G4_mul2_G16_mul0_G256_inv0 & m1_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p3_comar1_G4_mul2_G16_mul0_G256_inv0 = (m3_comar1_G4_mul2_G16_mul0_G256_inv0 & m2_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p1_comar1_G4_mul2_G16_mul0_G256_inv0 = (m0_comar1_G4_mul2_G16_mul0_G256_inv0 & m2_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p4_comar1_G4_mul2_G16_mul0_G256_inv0 = (m3_comar1_G4_mul2_G16_mul0_G256_inv0 & m1_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i0_comar1_G4_mul2_G16_mul0_G256_inv0 = (p1_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i1_comar1_G4_mul2_G16_mul0_G256_inv0 = (p2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i2_comar1_G4_mul2_G16_mul0_G256_inv0 = (p3_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i3_comar1_G4_mul2_G16_mul0_G256_inv0 = (p4_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0 = (i1_comar1_G4_mul2_G16_mul0_G256_inv0 ^ i2_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0 = (i0_comar1_G4_mul2_G16_mul0_G256_inv0 ^ i3_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p0_0_G4_mul2_G16_mul0_G256_inv0 = (i1xori2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_1_comar1_G4_mul2_G16_mul0_G256_inv0 = (r00_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p1_0_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul0_G256_inv0);
    assign p0_G4_mul2_G16_mul0_G256_inv0 = (p0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign p1_G4_mul2_G16_mul0_G256_inv0 = (p1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul0_G256_inv0 = (r00_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r10_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r20_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r30_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r40_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul0_G256_inv0 = (r50_G4_mul2_G16_mul0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul0_G256_inv0 = (b0_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul0_G256_inv0 = (d1_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul0_G256_inv0 = (d0_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign m3_comar2_G4_mul2_G16_mul0_G256_inv0 = (b1_G4_mul2_G16_mul0_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign p2_comar2_G4_mul2_G16_mul0_G256_inv0 = (m0_comar2_G4_mul2_G16_mul0_G256_inv0 & m1_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign p3_comar2_G4_mul2_G16_mul0_G256_inv0 = (m3_comar2_G4_mul2_G16_mul0_G256_inv0 & m2_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign p1_comar2_G4_mul2_G16_mul0_G256_inv0 = (m0_comar2_G4_mul2_G16_mul0_G256_inv0 & m2_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign p4_comar2_G4_mul2_G16_mul0_G256_inv0 = (m3_comar2_G4_mul2_G16_mul0_G256_inv0 & m1_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i0_comar2_G4_mul2_G16_mul0_G256_inv0 = (p1_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i1_comar2_G4_mul2_G16_mul0_G256_inv0 = (p2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i2_comar2_G4_mul2_G16_mul0_G256_inv0 = (p3_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i3_comar2_G4_mul2_G16_mul0_G256_inv0 = (p4_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0 = (i1_comar2_G4_mul2_G16_mul0_G256_inv0 ^ i2_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0 = (i0_comar2_G4_mul2_G16_mul0_G256_inv0 ^ i3_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign q0_0_G4_mul2_G16_mul0_G256_inv0 = (i1xori2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_1_comar2_G4_mul2_G16_mul0_G256_inv0 = (r00_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul0_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G4_mul2_G16_mul0_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul0_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G4_mul2_G16_mul0_G256_inv0 = (q0_0_G4_mul2_G16_mul0_G256_inv0 ^ e0_G4_mul2_G16_mul0_G256_inv0);
    assign q1_G4_mul2_G16_mul0_G256_inv0 = (q1_0_G4_mul2_G16_mul0_G256_inv0 ^ e1_G4_mul2_G16_mul0_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul0_G256_inv0 = (p1_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul2_G16_mul0_G256_inv0 = (p0_G4_mul2_G16_mul0_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul0_G256_inv0 = (p1ls1_G4_mul2_G16_mul0_G256_inv0 | q1_G4_mul2_G16_mul0_G256_inv0);
    assign q1_0_G16_mul0_G256_inv0 = (p0ls1_G4_mul2_G16_mul0_G256_inv0 | q0_G4_mul2_G16_mul0_G256_inv0);
    assign q0_G16_mul0_G256_inv0 = (q0_0_G16_mul0_G256_inv0 ^ e01_G16_mul0_G256_inv0);
    assign q1_G16_mul0_G256_inv0 = (q1_0_G16_mul0_G256_inv0 ^ e11_G16_mul0_G256_inv0);
    assign p0ls2_G16_mul0_G256_inv0 = (p0_G16_mul0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_mul0_G256_inv0 = (p1_G16_mul0_G256_inv0 << dec_2_inp);
    assign d0_G256_inv0 = (p0ls2_G16_mul0_G256_inv0 | q0_G16_mul0_G256_inv0);
    assign d1_G256_inv0 = (p1ls2_G16_mul0_G256_inv0 | q1_G16_mul0_G256_inv0);
    assign c0xord0_G256_inv0 = (c0_G256_inv0 ^ d0_G256_inv0);
    assign c1xord1_G256_inv0 = (c1_G256_inv0 ^ d1_G256_inv0);
    assign r00_G16_inv0_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_inv0_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_inv0_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_inv0_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_inv0_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_inv0_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & dec_12_inp);
    assign a0_G16_inv0_G256_inv0 = (a0_0_G16_inv0_G256_inv0 >> dec_2_inp);
    assign a1_G16_inv0_G256_inv0 = (a1_0_G16_inv0_G256_inv0 >> dec_2_inp);
    assign b0_G16_inv0_G256_inv0 = (c0xord0_G256_inv0 & dec_3_inp);
    assign b1_G16_inv0_G256_inv0 = (c1xord1_G256_inv0 & dec_3_inp);
    assign a0xorb0_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 ^ b0_G16_inv0_G256_inv0);
    assign a1xorb1_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 ^ b1_G16_inv0_G256_inv0);
    assign a0_0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq2_G16_inv0_G256_inv0 = (a0_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq2_G16_inv0_G256_inv0 = (a1_0_G4_sq2_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq2_G16_inv0_G256_inv0 = (a0xorb0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq2_G16_inv0_G256_inv0 = (a1xorb1_G16_inv0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq2_G16_inv0_G256_inv0 = (b0_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq2_G16_inv0_G256_inv0 = (b1_G4_sq2_G16_inv0_G256_inv0 << dec_1_inp);
    assign c0_0_G16_inv0_G256_inv0 = (b0ls1_G4_sq2_G16_inv0_G256_inv0 | a0_G4_sq2_G16_inv0_G256_inv0);
    assign c1_0_G16_inv0_G256_inv0 = (b1ls1_G4_sq2_G16_inv0_G256_inv0 | a1_G4_sq2_G16_inv0_G256_inv0);
    assign a0_0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_0_G4_scl_N1_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N1_G16_inv0_G256_inv0 = (c0_0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N1_G16_inv0_G256_inv0 = (c1_0_G16_inv0_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N1_G16_inv0_G256_inv0 = b0_G4_scl_N1_G16_inv0_G256_inv0;
    assign p1_G4_scl_N1_G16_inv0_G256_inv0 = b1_G4_scl_N1_G16_inv0_G256_inv0;
    assign q0_G4_scl_N1_G16_inv0_G256_inv0 = (a0_G4_scl_N1_G16_inv0_G256_inv0 ^ b0_G4_scl_N1_G16_inv0_G256_inv0);
    assign q1_G4_scl_N1_G16_inv0_G256_inv0 = (a1_G4_scl_N1_G16_inv0_G256_inv0 ^ b1_G4_scl_N1_G16_inv0_G256_inv0);
    assign p1ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p1_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N1_G16_inv0_G256_inv0 = (p0_G4_scl_N1_G16_inv0_G256_inv0 << dec_1_inp);
    assign c0_G16_inv0_G256_inv0 = (p0ls1_G4_scl_N1_G16_inv0_G256_inv0 | q0_G4_scl_N1_G16_inv0_G256_inv0);
    assign c1_G16_inv0_G256_inv0 = (p1ls1_G4_scl_N1_G16_inv0_G256_inv0 | q1_G4_scl_N1_G16_inv0_G256_inv0);
    assign r00_G4_mul3_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul3_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul3_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul3_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul3_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul3_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul3_G16_inv0_G256_inv0 = (a0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul3_G16_inv0_G256_inv0 = (a1_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul3_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul3_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul3_G16_inv0_G256_inv0 = (c0_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul3_G16_inv0_G256_inv0 = (c1_0_G4_mul3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul3_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul3_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ b0_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ d0_G4_mul3_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ b1_G4_mul3_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ d1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul3_G16_inv0_G256_inv0 = (axorb_0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign m1_comar0_G4_mul3_G16_inv0_G256_inv0 = (cxord_1_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign m2_comar0_G4_mul3_G16_inv0_G256_inv0 = (cxord_0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign m3_comar0_G4_mul3_G16_inv0_G256_inv0 = (axorb_1_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign p2_comar0_G4_mul3_G16_inv0_G256_inv0 = (m0_comar0_G4_mul3_G16_inv0_G256_inv0 & m1_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign p3_comar0_G4_mul3_G16_inv0_G256_inv0 = (m3_comar0_G4_mul3_G16_inv0_G256_inv0 & m2_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_comar0_G4_mul3_G16_inv0_G256_inv0 = (m0_comar0_G4_mul3_G16_inv0_G256_inv0 & m2_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign p4_comar0_G4_mul3_G16_inv0_G256_inv0 = (m3_comar0_G4_mul3_G16_inv0_G256_inv0 & m1_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i0_comar0_G4_mul3_G16_inv0_G256_inv0 = (p1_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i1_comar0_G4_mul3_G16_inv0_G256_inv0 = (p2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i2_comar0_G4_mul3_G16_inv0_G256_inv0 = (p3_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i3_comar0_G4_mul3_G16_inv0_G256_inv0 = (p4_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0 = (i1_comar0_G4_mul3_G16_inv0_G256_inv0 ^ i2_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0 = (i0_comar0_G4_mul3_G16_inv0_G256_inv0 ^ i3_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign e0_G4_mul3_G16_inv0_G256_inv0 = (i1xori2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_1_comar0_G4_mul3_G16_inv0_G256_inv0 = (r00_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign e1_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul3_G16_inv0_G256_inv0 = (a0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign m1_comar1_G4_mul3_G16_inv0_G256_inv0 = (c1_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign m2_comar1_G4_mul3_G16_inv0_G256_inv0 = (c0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign m3_comar1_G4_mul3_G16_inv0_G256_inv0 = (a1_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p2_comar1_G4_mul3_G16_inv0_G256_inv0 = (m0_comar1_G4_mul3_G16_inv0_G256_inv0 & m1_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p3_comar1_G4_mul3_G16_inv0_G256_inv0 = (m3_comar1_G4_mul3_G16_inv0_G256_inv0 & m2_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p1_comar1_G4_mul3_G16_inv0_G256_inv0 = (m0_comar1_G4_mul3_G16_inv0_G256_inv0 & m2_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p4_comar1_G4_mul3_G16_inv0_G256_inv0 = (m3_comar1_G4_mul3_G16_inv0_G256_inv0 & m1_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i0_comar1_G4_mul3_G16_inv0_G256_inv0 = (p1_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i1_comar1_G4_mul3_G16_inv0_G256_inv0 = (p2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i2_comar1_G4_mul3_G16_inv0_G256_inv0 = (p3_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i3_comar1_G4_mul3_G16_inv0_G256_inv0 = (p4_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0 = (i1_comar1_G4_mul3_G16_inv0_G256_inv0 ^ i2_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0 = (i0_comar1_G4_mul3_G16_inv0_G256_inv0 ^ i3_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p0_0_G4_mul3_G16_inv0_G256_inv0 = (i1xori2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_1_comar1_G4_mul3_G16_inv0_G256_inv0 = (r00_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p1_0_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul3_G16_inv0_G256_inv0);
    assign p0_G4_mul3_G16_inv0_G256_inv0 = (p0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign p1_G4_mul3_G16_inv0_G256_inv0 = (p1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul3_G16_inv0_G256_inv0 = (r00_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r10_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r20_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r30_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r40_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul3_G16_inv0_G256_inv0 = (r50_G4_mul3_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul3_G16_inv0_G256_inv0 = (b0_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign m1_comar2_G4_mul3_G16_inv0_G256_inv0 = (d1_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign m2_comar2_G4_mul3_G16_inv0_G256_inv0 = (d0_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign m3_comar2_G4_mul3_G16_inv0_G256_inv0 = (b1_G4_mul3_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign p2_comar2_G4_mul3_G16_inv0_G256_inv0 = (m0_comar2_G4_mul3_G16_inv0_G256_inv0 & m1_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign p3_comar2_G4_mul3_G16_inv0_G256_inv0 = (m3_comar2_G4_mul3_G16_inv0_G256_inv0 & m2_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign p1_comar2_G4_mul3_G16_inv0_G256_inv0 = (m0_comar2_G4_mul3_G16_inv0_G256_inv0 & m2_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign p4_comar2_G4_mul3_G16_inv0_G256_inv0 = (m3_comar2_G4_mul3_G16_inv0_G256_inv0 & m1_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i0_comar2_G4_mul3_G16_inv0_G256_inv0 = (p1_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i1_comar2_G4_mul3_G16_inv0_G256_inv0 = (p2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i2_comar2_G4_mul3_G16_inv0_G256_inv0 = (p3_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i3_comar2_G4_mul3_G16_inv0_G256_inv0 = (p4_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0 = (i1_comar2_G4_mul3_G16_inv0_G256_inv0 ^ i2_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0 = (i0_comar2_G4_mul3_G16_inv0_G256_inv0 ^ i3_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign q0_0_G4_mul3_G16_inv0_G256_inv0 = (i1xori2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_1_comar2_G4_mul3_G16_inv0_G256_inv0 = (r00_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul3_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign q1_0_G4_mul3_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul3_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul3_G16_inv0_G256_inv0);
    assign q0_G4_mul3_G16_inv0_G256_inv0 = (q0_0_G4_mul3_G16_inv0_G256_inv0 ^ e0_G4_mul3_G16_inv0_G256_inv0);
    assign q1_G4_mul3_G16_inv0_G256_inv0 = (q1_0_G4_mul3_G16_inv0_G256_inv0 ^ e1_G4_mul3_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul3_G16_inv0_G256_inv0 = (p1_G4_mul3_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul3_G16_inv0_G256_inv0 = (p0_G4_mul3_G16_inv0_G256_inv0 << dec_1_inp);
    assign d0_G16_inv0_G256_inv0 = (p1ls1_G4_mul3_G16_inv0_G256_inv0 | q1_G4_mul3_G16_inv0_G256_inv0);
    assign d1_G16_inv0_G256_inv0 = (p0ls1_G4_mul3_G16_inv0_G256_inv0 | q0_G4_mul3_G16_inv0_G256_inv0);
    assign c0xord0_G16_inv0_G256_inv0 = (c0_G16_inv0_G256_inv0 ^ d0_G16_inv0_G256_inv0);
    assign c1xord1_G16_inv0_G256_inv0 = (c1_G16_inv0_G256_inv0 ^ d1_G16_inv0_G256_inv0);
    assign a0_0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_sq3_G16_inv0_G256_inv0 = (a0_0_G4_sq3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_sq3_G16_inv0_G256_inv0 = (a1_0_G4_sq3_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_sq3_G16_inv0_G256_inv0 = (c0xord0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_sq3_G16_inv0_G256_inv0 = (c1xord1_G16_inv0_G256_inv0 & dec_1_inp);
    assign b0ls1_G4_sq3_G16_inv0_G256_inv0 = (b0_G4_sq3_G16_inv0_G256_inv0 << dec_1_inp);
    assign b1ls1_G4_sq3_G16_inv0_G256_inv0 = (b1_G4_sq3_G16_inv0_G256_inv0 << dec_1_inp);
    assign e0_G16_inv0_G256_inv0 = (b0ls1_G4_sq3_G16_inv0_G256_inv0 | a0_G4_sq3_G16_inv0_G256_inv0);
    assign e1_G16_inv0_G256_inv0 = (b1ls1_G4_sq3_G16_inv0_G256_inv0 | a1_G4_sq3_G16_inv0_G256_inv0);
    assign r00_G4_mul4_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul4_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul4_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul4_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul4_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul4_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul4_G16_inv0_G256_inv0 = (a0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul4_G16_inv0_G256_inv0 = (a1_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul4_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul4_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul4_G16_inv0_G256_inv0 = (c0_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul4_G16_inv0_G256_inv0 = (c1_0_G4_mul4_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul4_G16_inv0_G256_inv0 = (b0_G16_inv0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul4_G16_inv0_G256_inv0 = (b1_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ b0_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ d0_G4_mul4_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ b1_G4_mul4_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ d1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul4_G16_inv0_G256_inv0 = (axorb_0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign m1_comar0_G4_mul4_G16_inv0_G256_inv0 = (cxord_1_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign m2_comar0_G4_mul4_G16_inv0_G256_inv0 = (cxord_0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign m3_comar0_G4_mul4_G16_inv0_G256_inv0 = (axorb_1_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign p2_comar0_G4_mul4_G16_inv0_G256_inv0 = (m0_comar0_G4_mul4_G16_inv0_G256_inv0 & m1_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign p3_comar0_G4_mul4_G16_inv0_G256_inv0 = (m3_comar0_G4_mul4_G16_inv0_G256_inv0 & m2_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_comar0_G4_mul4_G16_inv0_G256_inv0 = (m0_comar0_G4_mul4_G16_inv0_G256_inv0 & m2_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign p4_comar0_G4_mul4_G16_inv0_G256_inv0 = (m3_comar0_G4_mul4_G16_inv0_G256_inv0 & m1_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i0_comar0_G4_mul4_G16_inv0_G256_inv0 = (p1_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i1_comar0_G4_mul4_G16_inv0_G256_inv0 = (p2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i2_comar0_G4_mul4_G16_inv0_G256_inv0 = (p3_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i3_comar0_G4_mul4_G16_inv0_G256_inv0 = (p4_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0 = (i1_comar0_G4_mul4_G16_inv0_G256_inv0 ^ i2_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0 = (i0_comar0_G4_mul4_G16_inv0_G256_inv0 ^ i3_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign e0_G4_mul4_G16_inv0_G256_inv0 = (i1xori2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_1_comar0_G4_mul4_G16_inv0_G256_inv0 = (r00_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign e1_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul4_G16_inv0_G256_inv0 = (a0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign m1_comar1_G4_mul4_G16_inv0_G256_inv0 = (c1_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign m2_comar1_G4_mul4_G16_inv0_G256_inv0 = (c0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign m3_comar1_G4_mul4_G16_inv0_G256_inv0 = (a1_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p2_comar1_G4_mul4_G16_inv0_G256_inv0 = (m0_comar1_G4_mul4_G16_inv0_G256_inv0 & m1_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p3_comar1_G4_mul4_G16_inv0_G256_inv0 = (m3_comar1_G4_mul4_G16_inv0_G256_inv0 & m2_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_comar1_G4_mul4_G16_inv0_G256_inv0 = (m0_comar1_G4_mul4_G16_inv0_G256_inv0 & m2_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p4_comar1_G4_mul4_G16_inv0_G256_inv0 = (m3_comar1_G4_mul4_G16_inv0_G256_inv0 & m1_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i0_comar1_G4_mul4_G16_inv0_G256_inv0 = (p1_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i1_comar1_G4_mul4_G16_inv0_G256_inv0 = (p2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i2_comar1_G4_mul4_G16_inv0_G256_inv0 = (p3_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i3_comar1_G4_mul4_G16_inv0_G256_inv0 = (p4_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0 = (i1_comar1_G4_mul4_G16_inv0_G256_inv0 ^ i2_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0 = (i0_comar1_G4_mul4_G16_inv0_G256_inv0 ^ i3_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p0_0_G4_mul4_G16_inv0_G256_inv0 = (i1xori2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_1_comar1_G4_mul4_G16_inv0_G256_inv0 = (r00_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_0_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul4_G16_inv0_G256_inv0);
    assign p0_G4_mul4_G16_inv0_G256_inv0 = (p0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G4_mul4_G16_inv0_G256_inv0 = (p1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul4_G16_inv0_G256_inv0 = (r00_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r10_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r20_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r30_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r40_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul4_G16_inv0_G256_inv0 = (r50_G4_mul4_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul4_G16_inv0_G256_inv0 = (b0_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign m1_comar2_G4_mul4_G16_inv0_G256_inv0 = (d1_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign m2_comar2_G4_mul4_G16_inv0_G256_inv0 = (d0_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign m3_comar2_G4_mul4_G16_inv0_G256_inv0 = (b1_G4_mul4_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign p2_comar2_G4_mul4_G16_inv0_G256_inv0 = (m0_comar2_G4_mul4_G16_inv0_G256_inv0 & m1_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign p3_comar2_G4_mul4_G16_inv0_G256_inv0 = (m3_comar2_G4_mul4_G16_inv0_G256_inv0 & m2_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign p1_comar2_G4_mul4_G16_inv0_G256_inv0 = (m0_comar2_G4_mul4_G16_inv0_G256_inv0 & m2_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign p4_comar2_G4_mul4_G16_inv0_G256_inv0 = (m3_comar2_G4_mul4_G16_inv0_G256_inv0 & m1_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i0_comar2_G4_mul4_G16_inv0_G256_inv0 = (p1_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i1_comar2_G4_mul4_G16_inv0_G256_inv0 = (p2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i2_comar2_G4_mul4_G16_inv0_G256_inv0 = (p3_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i3_comar2_G4_mul4_G16_inv0_G256_inv0 = (p4_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0 = (i1_comar2_G4_mul4_G16_inv0_G256_inv0 ^ i2_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0 = (i0_comar2_G4_mul4_G16_inv0_G256_inv0 ^ i3_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign q0_0_G4_mul4_G16_inv0_G256_inv0 = (i1xori2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_1_comar2_G4_mul4_G16_inv0_G256_inv0 = (r00_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul4_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign q1_0_G4_mul4_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul4_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul4_G16_inv0_G256_inv0);
    assign q0_G4_mul4_G16_inv0_G256_inv0 = (q0_0_G4_mul4_G16_inv0_G256_inv0 ^ e0_G4_mul4_G16_inv0_G256_inv0);
    assign q1_G4_mul4_G16_inv0_G256_inv0 = (q1_0_G4_mul4_G16_inv0_G256_inv0 ^ e1_G4_mul4_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul4_G16_inv0_G256_inv0 = (p1_G4_mul4_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul4_G16_inv0_G256_inv0 = (p0_G4_mul4_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0_G16_inv0_G256_inv0 = (p1ls1_G4_mul4_G16_inv0_G256_inv0 | q1_G4_mul4_G16_inv0_G256_inv0);
    assign p1_G16_inv0_G256_inv0 = (p0ls1_G4_mul4_G16_inv0_G256_inv0 | q0_G4_mul4_G16_inv0_G256_inv0);
    assign r00_G4_mul5_G16_inv0_G256_inv0 = (r00_G16_inv0_G256_inv0 % dec_4_inp);
    assign r10_G4_mul5_G16_inv0_G256_inv0 = (r10_G16_inv0_G256_inv0 % dec_4_inp);
    assign r20_G4_mul5_G16_inv0_G256_inv0 = (r20_G16_inv0_G256_inv0 % dec_4_inp);
    assign r30_G4_mul5_G16_inv0_G256_inv0 = (r30_G16_inv0_G256_inv0 % dec_4_inp);
    assign r40_G4_mul5_G16_inv0_G256_inv0 = (r40_G16_inv0_G256_inv0 % dec_4_inp);
    assign r50_G4_mul5_G16_inv0_G256_inv0 = (r50_G16_inv0_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & dec_2_inp);
    assign a0_G4_mul5_G16_inv0_G256_inv0 = (a0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul5_G16_inv0_G256_inv0 = (a1_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul5_G16_inv0_G256_inv0 = (e0_G16_inv0_G256_inv0 & dec_1_inp);
    assign b1_G4_mul5_G16_inv0_G256_inv0 = (e1_G16_inv0_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_2_inp);
    assign c0_G4_mul5_G16_inv0_G256_inv0 = (c0_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul5_G16_inv0_G256_inv0 = (c1_0_G4_mul5_G16_inv0_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul5_G16_inv0_G256_inv0 = (a0_G16_inv0_G256_inv0 & dec_1_inp);
    assign d1_G4_mul5_G16_inv0_G256_inv0 = (a1_G16_inv0_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ b0_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_0_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ d0_G4_mul5_G16_inv0_G256_inv0);
    assign axorb_1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ b1_G4_mul5_G16_inv0_G256_inv0);
    assign cxord_1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ d1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar0_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul5_G16_inv0_G256_inv0 = (axorb_0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign m1_comar0_G4_mul5_G16_inv0_G256_inv0 = (cxord_1_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign m2_comar0_G4_mul5_G16_inv0_G256_inv0 = (cxord_0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign m3_comar0_G4_mul5_G16_inv0_G256_inv0 = (axorb_1_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign p2_comar0_G4_mul5_G16_inv0_G256_inv0 = (m0_comar0_G4_mul5_G16_inv0_G256_inv0 & m1_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign p3_comar0_G4_mul5_G16_inv0_G256_inv0 = (m3_comar0_G4_mul5_G16_inv0_G256_inv0 & m2_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_comar0_G4_mul5_G16_inv0_G256_inv0 = (m0_comar0_G4_mul5_G16_inv0_G256_inv0 & m2_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign p4_comar0_G4_mul5_G16_inv0_G256_inv0 = (m3_comar0_G4_mul5_G16_inv0_G256_inv0 & m1_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i0_comar0_G4_mul5_G16_inv0_G256_inv0 = (p1_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i1_comar0_G4_mul5_G16_inv0_G256_inv0 = (p2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i2_comar0_G4_mul5_G16_inv0_G256_inv0 = (p3_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i3_comar0_G4_mul5_G16_inv0_G256_inv0 = (p4_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0 = (i1_comar0_G4_mul5_G16_inv0_G256_inv0 ^ i2_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0 = (i0_comar0_G4_mul5_G16_inv0_G256_inv0 ^ i3_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign e0_G4_mul5_G16_inv0_G256_inv0 = (i1xori2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_1_comar0_G4_mul5_G16_inv0_G256_inv0 = (r00_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar0_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign e1_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar0_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar0_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar1_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul5_G16_inv0_G256_inv0 = (a0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign m1_comar1_G4_mul5_G16_inv0_G256_inv0 = (c1_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign m2_comar1_G4_mul5_G16_inv0_G256_inv0 = (c0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign m3_comar1_G4_mul5_G16_inv0_G256_inv0 = (a1_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p2_comar1_G4_mul5_G16_inv0_G256_inv0 = (m0_comar1_G4_mul5_G16_inv0_G256_inv0 & m1_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p3_comar1_G4_mul5_G16_inv0_G256_inv0 = (m3_comar1_G4_mul5_G16_inv0_G256_inv0 & m2_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p1_comar1_G4_mul5_G16_inv0_G256_inv0 = (m0_comar1_G4_mul5_G16_inv0_G256_inv0 & m2_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p4_comar1_G4_mul5_G16_inv0_G256_inv0 = (m3_comar1_G4_mul5_G16_inv0_G256_inv0 & m1_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i0_comar1_G4_mul5_G16_inv0_G256_inv0 = (p1_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i1_comar1_G4_mul5_G16_inv0_G256_inv0 = (p2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i2_comar1_G4_mul5_G16_inv0_G256_inv0 = (p3_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i3_comar1_G4_mul5_G16_inv0_G256_inv0 = (p4_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0 = (i1_comar1_G4_mul5_G16_inv0_G256_inv0 ^ i2_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0 = (i0_comar1_G4_mul5_G16_inv0_G256_inv0 ^ i3_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p0_0_G4_mul5_G16_inv0_G256_inv0 = (i1xori2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_1_comar1_G4_mul5_G16_inv0_G256_inv0 = (r00_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar1_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p1_0_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar1_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar1_G4_mul5_G16_inv0_G256_inv0);
    assign p0_G4_mul5_G16_inv0_G256_inv0 = (p0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign p1_G4_mul5_G16_inv0_G256_inv0 = (p1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign r00_comar2_G4_mul5_G16_inv0_G256_inv0 = (r00_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r10_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r20_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r30_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r40_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul5_G16_inv0_G256_inv0 = (r50_G4_mul5_G16_inv0_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul5_G16_inv0_G256_inv0 = (b0_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign m1_comar2_G4_mul5_G16_inv0_G256_inv0 = (d1_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign m2_comar2_G4_mul5_G16_inv0_G256_inv0 = (d0_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign m3_comar2_G4_mul5_G16_inv0_G256_inv0 = (b1_G4_mul5_G16_inv0_G256_inv0 ^ r00_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign p2_comar2_G4_mul5_G16_inv0_G256_inv0 = (m0_comar2_G4_mul5_G16_inv0_G256_inv0 & m1_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign p3_comar2_G4_mul5_G16_inv0_G256_inv0 = (m3_comar2_G4_mul5_G16_inv0_G256_inv0 & m2_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign p1_comar2_G4_mul5_G16_inv0_G256_inv0 = (m0_comar2_G4_mul5_G16_inv0_G256_inv0 & m2_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign p4_comar2_G4_mul5_G16_inv0_G256_inv0 = (m3_comar2_G4_mul5_G16_inv0_G256_inv0 & m1_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i0_comar2_G4_mul5_G16_inv0_G256_inv0 = (p1_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i1_comar2_G4_mul5_G16_inv0_G256_inv0 = (p2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i2_comar2_G4_mul5_G16_inv0_G256_inv0 = (p3_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i3_comar2_G4_mul5_G16_inv0_G256_inv0 = (p4_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0 = (i1_comar2_G4_mul5_G16_inv0_G256_inv0 ^ i2_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0 = (i0_comar2_G4_mul5_G16_inv0_G256_inv0 ^ i3_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign q0_0_G4_mul5_G16_inv0_G256_inv0 = (i1xori2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ i0xori3_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_1_comar2_G4_mul5_G16_inv0_G256_inv0 = (r00_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_2_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_1_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r0_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_3_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_2_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r1_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign y1_4_comar2_G4_mul5_G16_inv0_G256_inv0 = (y1_3_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r2_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign q1_0_G4_mul5_G16_inv0_G256_inv0 = (y1_4_comar2_G4_mul5_G16_inv0_G256_inv0 ^ r3_10_comar2_G4_mul5_G16_inv0_G256_inv0);
    assign q0_G4_mul5_G16_inv0_G256_inv0 = (q0_0_G4_mul5_G16_inv0_G256_inv0 ^ e0_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G4_mul5_G16_inv0_G256_inv0 = (q1_0_G4_mul5_G16_inv0_G256_inv0 ^ e1_G4_mul5_G16_inv0_G256_inv0);
    assign p1ls1_G4_mul5_G16_inv0_G256_inv0 = (p1_G4_mul5_G16_inv0_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul5_G16_inv0_G256_inv0 = (p0_G4_mul5_G16_inv0_G256_inv0 << dec_1_inp);
    assign q0_G16_inv0_G256_inv0 = (p1ls1_G4_mul5_G16_inv0_G256_inv0 | q1_G4_mul5_G16_inv0_G256_inv0);
    assign q1_G16_inv0_G256_inv0 = (p0ls1_G4_mul5_G16_inv0_G256_inv0 | q0_G4_mul5_G16_inv0_G256_inv0);
    assign p0ls2_G16_inv0_G256_inv0 = (p0_G16_inv0_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_inv0_G256_inv0 = (p1_G16_inv0_G256_inv0 << dec_2_inp);
    assign e0_G256_inv0 = (p0ls2_G16_inv0_G256_inv0 | q0_G16_inv0_G256_inv0);
    assign e1_G256_inv0 = (p1ls2_G16_inv0_G256_inv0 | q1_G16_inv0_G256_inv0);
    assign r00_G16_mul1_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul1_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul1_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul1_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul1_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul1_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul1_G256_inv0 = (e1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul1_G256_inv0 = (a0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul1_G256_inv0 = (a1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul1_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul1_G256_inv0 = (e1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul1_G256_inv0 = (c0_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul1_G256_inv0 = (c1_0_G16_mul1_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul1_G256_inv0 = (b0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul1_G256_inv0 = (b1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 ^ b0_G16_mul1_G256_inv0);
    assign cxord_0_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 ^ d0_G16_mul1_G256_inv0);
    assign axorb_1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 ^ b1_G16_mul1_G256_inv0);
    assign cxord_1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 ^ d1_G16_mul1_G256_inv0);
    assign r00_G4_mul0_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul1_G256_inv0 = (a0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul1_G256_inv0 = (a1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul1_G256_inv0 = (c0_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul1_G256_inv0 = (c1_0_G4_mul0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ b0_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ d0_G4_mul0_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ b1_G4_mul0_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ d1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul1_G256_inv0 = (axorb_0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul1_G256_inv0 = (cxord_1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul1_G256_inv0 = (cxord_0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign m3_comar0_G4_mul0_G16_mul1_G256_inv0 = (axorb_1_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign p2_comar0_G4_mul0_G16_mul1_G256_inv0 = (m0_comar0_G4_mul0_G16_mul1_G256_inv0 & m1_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign p3_comar0_G4_mul0_G16_mul1_G256_inv0 = (m3_comar0_G4_mul0_G16_mul1_G256_inv0 & m2_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_comar0_G4_mul0_G16_mul1_G256_inv0 = (m0_comar0_G4_mul0_G16_mul1_G256_inv0 & m2_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign p4_comar0_G4_mul0_G16_mul1_G256_inv0 = (m3_comar0_G4_mul0_G16_mul1_G256_inv0 & m1_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i0_comar0_G4_mul0_G16_mul1_G256_inv0 = (p1_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i1_comar0_G4_mul0_G16_mul1_G256_inv0 = (p2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i2_comar0_G4_mul0_G16_mul1_G256_inv0 = (p3_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i3_comar0_G4_mul0_G16_mul1_G256_inv0 = (p4_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0 = (i1_comar0_G4_mul0_G16_mul1_G256_inv0 ^ i2_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0 = (i0_comar0_G4_mul0_G16_mul1_G256_inv0 ^ i3_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign e0_G4_mul0_G16_mul1_G256_inv0 = (i1xori2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_1_comar0_G4_mul0_G16_mul1_G256_inv0 = (r00_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul1_G256_inv0 = (a0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul1_G256_inv0 = (c1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul1_G256_inv0 = (c0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign m3_comar1_G4_mul0_G16_mul1_G256_inv0 = (a1_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p2_comar1_G4_mul0_G16_mul1_G256_inv0 = (m0_comar1_G4_mul0_G16_mul1_G256_inv0 & m1_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p3_comar1_G4_mul0_G16_mul1_G256_inv0 = (m3_comar1_G4_mul0_G16_mul1_G256_inv0 & m2_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p1_comar1_G4_mul0_G16_mul1_G256_inv0 = (m0_comar1_G4_mul0_G16_mul1_G256_inv0 & m2_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p4_comar1_G4_mul0_G16_mul1_G256_inv0 = (m3_comar1_G4_mul0_G16_mul1_G256_inv0 & m1_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i0_comar1_G4_mul0_G16_mul1_G256_inv0 = (p1_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i1_comar1_G4_mul0_G16_mul1_G256_inv0 = (p2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i2_comar1_G4_mul0_G16_mul1_G256_inv0 = (p3_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i3_comar1_G4_mul0_G16_mul1_G256_inv0 = (p4_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0 = (i1_comar1_G4_mul0_G16_mul1_G256_inv0 ^ i2_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0 = (i0_comar1_G4_mul0_G16_mul1_G256_inv0 ^ i3_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p0_0_G4_mul0_G16_mul1_G256_inv0 = (i1xori2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_1_comar1_G4_mul0_G16_mul1_G256_inv0 = (r00_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p1_0_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul1_G256_inv0);
    assign p0_G4_mul0_G16_mul1_G256_inv0 = (p0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign p1_G4_mul0_G16_mul1_G256_inv0 = (p1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul1_G256_inv0 = (r00_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r10_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r20_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r30_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r40_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul1_G256_inv0 = (r50_G4_mul0_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul1_G256_inv0 = (b0_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul1_G256_inv0 = (d1_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul1_G256_inv0 = (d0_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign m3_comar2_G4_mul0_G16_mul1_G256_inv0 = (b1_G4_mul0_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign p2_comar2_G4_mul0_G16_mul1_G256_inv0 = (m0_comar2_G4_mul0_G16_mul1_G256_inv0 & m1_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign p3_comar2_G4_mul0_G16_mul1_G256_inv0 = (m3_comar2_G4_mul0_G16_mul1_G256_inv0 & m2_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign p1_comar2_G4_mul0_G16_mul1_G256_inv0 = (m0_comar2_G4_mul0_G16_mul1_G256_inv0 & m2_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign p4_comar2_G4_mul0_G16_mul1_G256_inv0 = (m3_comar2_G4_mul0_G16_mul1_G256_inv0 & m1_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i0_comar2_G4_mul0_G16_mul1_G256_inv0 = (p1_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i1_comar2_G4_mul0_G16_mul1_G256_inv0 = (p2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i2_comar2_G4_mul0_G16_mul1_G256_inv0 = (p3_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i3_comar2_G4_mul0_G16_mul1_G256_inv0 = (p4_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0 = (i1_comar2_G4_mul0_G16_mul1_G256_inv0 ^ i2_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0 = (i0_comar2_G4_mul0_G16_mul1_G256_inv0 ^ i3_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign q0_0_G4_mul0_G16_mul1_G256_inv0 = (i1xori2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_1_comar2_G4_mul0_G16_mul1_G256_inv0 = (r00_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign q1_0_G4_mul0_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul1_G256_inv0);
    assign q0_G4_mul0_G16_mul1_G256_inv0 = (q0_0_G4_mul0_G16_mul1_G256_inv0 ^ e0_G4_mul0_G16_mul1_G256_inv0);
    assign q1_G4_mul0_G16_mul1_G256_inv0 = (q1_0_G4_mul0_G16_mul1_G256_inv0 ^ e1_G4_mul0_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul1_G256_inv0 = (p1_G4_mul0_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul0_G16_mul1_G256_inv0 = (p0_G4_mul0_G16_mul1_G256_inv0 << dec_1_inp);
    assign e0_G16_mul1_G256_inv0 = (p1ls1_G4_mul0_G16_mul1_G256_inv0 | q1_G4_mul0_G16_mul1_G256_inv0);
    assign e1_G16_mul1_G256_inv0 = (p0ls1_G4_mul0_G16_mul1_G256_inv0 | q0_G4_mul0_G16_mul1_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_0_G4_scl_N0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_0_G4_scl_N0_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul1_G256_inv0 = (e0_G16_mul1_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N0_G16_mul1_G256_inv0 = (e1_G16_mul1_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul1_G256_inv0 = b0_G4_scl_N0_G16_mul1_G256_inv0;
    assign p1_G4_scl_N0_G16_mul1_G256_inv0 = b1_G4_scl_N0_G16_mul1_G256_inv0;
    assign q0_G4_scl_N0_G16_mul1_G256_inv0 = (a0_G4_scl_N0_G16_mul1_G256_inv0 ^ b0_G4_scl_N0_G16_mul1_G256_inv0);
    assign q1_G4_scl_N0_G16_mul1_G256_inv0 = (a1_G4_scl_N0_G16_mul1_G256_inv0 ^ b1_G4_scl_N0_G16_mul1_G256_inv0);
    assign p1ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p1_G4_scl_N0_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N0_G16_mul1_G256_inv0 = (p0_G4_scl_N0_G16_mul1_G256_inv0 << dec_1_inp);
    assign e01_G16_mul1_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul1_G256_inv0 | q0_G4_scl_N0_G16_mul1_G256_inv0);
    assign e11_G16_mul1_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul1_G256_inv0 | q1_G4_scl_N0_G16_mul1_G256_inv0);
    assign r00_G4_mul1_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul1_G256_inv0 = (a0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul1_G256_inv0 = (a1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul1_G256_inv0 = (a0_G16_mul1_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul1_G256_inv0 = (a1_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul1_G256_inv0 = (c0_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul1_G256_inv0 = (c1_0_G4_mul1_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul1_G256_inv0 = (c0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul1_G256_inv0 = (c1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ b0_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ d0_G4_mul1_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ b1_G4_mul1_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ d1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul1_G256_inv0 = (axorb_0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul1_G256_inv0 = (cxord_1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul1_G256_inv0 = (cxord_0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign m3_comar0_G4_mul1_G16_mul1_G256_inv0 = (axorb_1_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign p2_comar0_G4_mul1_G16_mul1_G256_inv0 = (m0_comar0_G4_mul1_G16_mul1_G256_inv0 & m1_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign p3_comar0_G4_mul1_G16_mul1_G256_inv0 = (m3_comar0_G4_mul1_G16_mul1_G256_inv0 & m2_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_comar0_G4_mul1_G16_mul1_G256_inv0 = (m0_comar0_G4_mul1_G16_mul1_G256_inv0 & m2_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign p4_comar0_G4_mul1_G16_mul1_G256_inv0 = (m3_comar0_G4_mul1_G16_mul1_G256_inv0 & m1_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i0_comar0_G4_mul1_G16_mul1_G256_inv0 = (p1_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i1_comar0_G4_mul1_G16_mul1_G256_inv0 = (p2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i2_comar0_G4_mul1_G16_mul1_G256_inv0 = (p3_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i3_comar0_G4_mul1_G16_mul1_G256_inv0 = (p4_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0 = (i1_comar0_G4_mul1_G16_mul1_G256_inv0 ^ i2_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0 = (i0_comar0_G4_mul1_G16_mul1_G256_inv0 ^ i3_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign e0_G4_mul1_G16_mul1_G256_inv0 = (i1xori2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_1_comar0_G4_mul1_G16_mul1_G256_inv0 = (r00_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign e1_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul1_G256_inv0 = (a0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul1_G256_inv0 = (c1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul1_G256_inv0 = (c0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign m3_comar1_G4_mul1_G16_mul1_G256_inv0 = (a1_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p2_comar1_G4_mul1_G16_mul1_G256_inv0 = (m0_comar1_G4_mul1_G16_mul1_G256_inv0 & m1_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p3_comar1_G4_mul1_G16_mul1_G256_inv0 = (m3_comar1_G4_mul1_G16_mul1_G256_inv0 & m2_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_comar1_G4_mul1_G16_mul1_G256_inv0 = (m0_comar1_G4_mul1_G16_mul1_G256_inv0 & m2_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p4_comar1_G4_mul1_G16_mul1_G256_inv0 = (m3_comar1_G4_mul1_G16_mul1_G256_inv0 & m1_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i0_comar1_G4_mul1_G16_mul1_G256_inv0 = (p1_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i1_comar1_G4_mul1_G16_mul1_G256_inv0 = (p2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i2_comar1_G4_mul1_G16_mul1_G256_inv0 = (p3_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i3_comar1_G4_mul1_G16_mul1_G256_inv0 = (p4_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0 = (i1_comar1_G4_mul1_G16_mul1_G256_inv0 ^ i2_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0 = (i0_comar1_G4_mul1_G16_mul1_G256_inv0 ^ i3_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p0_0_G4_mul1_G16_mul1_G256_inv0 = (i1xori2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_1_comar1_G4_mul1_G16_mul1_G256_inv0 = (r00_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G4_mul1_G16_mul1_G256_inv0 = (p0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign p1_G4_mul1_G16_mul1_G256_inv0 = (p1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul1_G256_inv0 = (r00_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r10_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r20_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r30_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r40_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul1_G256_inv0 = (r50_G4_mul1_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul1_G256_inv0 = (b0_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul1_G256_inv0 = (d1_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul1_G256_inv0 = (d0_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign m3_comar2_G4_mul1_G16_mul1_G256_inv0 = (b1_G4_mul1_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign p2_comar2_G4_mul1_G16_mul1_G256_inv0 = (m0_comar2_G4_mul1_G16_mul1_G256_inv0 & m1_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign p3_comar2_G4_mul1_G16_mul1_G256_inv0 = (m3_comar2_G4_mul1_G16_mul1_G256_inv0 & m2_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign p1_comar2_G4_mul1_G16_mul1_G256_inv0 = (m0_comar2_G4_mul1_G16_mul1_G256_inv0 & m2_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign p4_comar2_G4_mul1_G16_mul1_G256_inv0 = (m3_comar2_G4_mul1_G16_mul1_G256_inv0 & m1_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i0_comar2_G4_mul1_G16_mul1_G256_inv0 = (p1_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i1_comar2_G4_mul1_G16_mul1_G256_inv0 = (p2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i2_comar2_G4_mul1_G16_mul1_G256_inv0 = (p3_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i3_comar2_G4_mul1_G16_mul1_G256_inv0 = (p4_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0 = (i1_comar2_G4_mul1_G16_mul1_G256_inv0 ^ i2_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0 = (i0_comar2_G4_mul1_G16_mul1_G256_inv0 ^ i3_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign q0_0_G4_mul1_G16_mul1_G256_inv0 = (i1xori2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_1_comar2_G4_mul1_G16_mul1_G256_inv0 = (r00_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign q1_0_G4_mul1_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul1_G256_inv0);
    assign q0_G4_mul1_G16_mul1_G256_inv0 = (q0_0_G4_mul1_G16_mul1_G256_inv0 ^ e0_G4_mul1_G16_mul1_G256_inv0);
    assign q1_G4_mul1_G16_mul1_G256_inv0 = (q1_0_G4_mul1_G16_mul1_G256_inv0 ^ e1_G4_mul1_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul1_G256_inv0 = (p1_G4_mul1_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul1_G16_mul1_G256_inv0 = (p0_G4_mul1_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul1_G16_mul1_G256_inv0 | q1_G4_mul1_G16_mul1_G256_inv0);
    assign p1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul1_G16_mul1_G256_inv0 | q0_G4_mul1_G16_mul1_G256_inv0);
    assign p0_G16_mul1_G256_inv0 = (p0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign p1_G16_mul1_G256_inv0 = (p1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign r00_G4_mul2_G16_mul1_G256_inv0 = (r00_G16_mul1_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul1_G256_inv0 = (r10_G16_mul1_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul1_G256_inv0 = (r20_G16_mul1_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul1_G256_inv0 = (r30_G16_mul1_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul1_G256_inv0 = (r40_G16_mul1_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul1_G256_inv0 = (r50_G16_mul1_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul1_G256_inv0 = (a0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul1_G256_inv0 = (a1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul1_G256_inv0 = (b0_G16_mul1_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul1_G256_inv0 = (b1_G16_mul1_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul1_G256_inv0 = (c0_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul1_G256_inv0 = (c1_0_G4_mul2_G16_mul1_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul1_G256_inv0 = (d0_G16_mul1_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul1_G256_inv0 = (d1_G16_mul1_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ b0_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ d0_G4_mul2_G16_mul1_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ b1_G4_mul2_G16_mul1_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ d1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul1_G256_inv0 = (axorb_0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul1_G256_inv0 = (cxord_1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul1_G256_inv0 = (cxord_0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign m3_comar0_G4_mul2_G16_mul1_G256_inv0 = (axorb_1_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign p2_comar0_G4_mul2_G16_mul1_G256_inv0 = (m0_comar0_G4_mul2_G16_mul1_G256_inv0 & m1_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign p3_comar0_G4_mul2_G16_mul1_G256_inv0 = (m3_comar0_G4_mul2_G16_mul1_G256_inv0 & m2_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_comar0_G4_mul2_G16_mul1_G256_inv0 = (m0_comar0_G4_mul2_G16_mul1_G256_inv0 & m2_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign p4_comar0_G4_mul2_G16_mul1_G256_inv0 = (m3_comar0_G4_mul2_G16_mul1_G256_inv0 & m1_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i0_comar0_G4_mul2_G16_mul1_G256_inv0 = (p1_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i1_comar0_G4_mul2_G16_mul1_G256_inv0 = (p2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i2_comar0_G4_mul2_G16_mul1_G256_inv0 = (p3_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i3_comar0_G4_mul2_G16_mul1_G256_inv0 = (p4_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0 = (i1_comar0_G4_mul2_G16_mul1_G256_inv0 ^ i2_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0 = (i0_comar0_G4_mul2_G16_mul1_G256_inv0 ^ i3_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign e0_G4_mul2_G16_mul1_G256_inv0 = (i1xori2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_1_comar0_G4_mul2_G16_mul1_G256_inv0 = (r00_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign e1_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul1_G256_inv0 = (a0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul1_G256_inv0 = (c1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul1_G256_inv0 = (c0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign m3_comar1_G4_mul2_G16_mul1_G256_inv0 = (a1_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p2_comar1_G4_mul2_G16_mul1_G256_inv0 = (m0_comar1_G4_mul2_G16_mul1_G256_inv0 & m1_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p3_comar1_G4_mul2_G16_mul1_G256_inv0 = (m3_comar1_G4_mul2_G16_mul1_G256_inv0 & m2_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p1_comar1_G4_mul2_G16_mul1_G256_inv0 = (m0_comar1_G4_mul2_G16_mul1_G256_inv0 & m2_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p4_comar1_G4_mul2_G16_mul1_G256_inv0 = (m3_comar1_G4_mul2_G16_mul1_G256_inv0 & m1_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i0_comar1_G4_mul2_G16_mul1_G256_inv0 = (p1_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i1_comar1_G4_mul2_G16_mul1_G256_inv0 = (p2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i2_comar1_G4_mul2_G16_mul1_G256_inv0 = (p3_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i3_comar1_G4_mul2_G16_mul1_G256_inv0 = (p4_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0 = (i1_comar1_G4_mul2_G16_mul1_G256_inv0 ^ i2_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0 = (i0_comar1_G4_mul2_G16_mul1_G256_inv0 ^ i3_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p0_0_G4_mul2_G16_mul1_G256_inv0 = (i1xori2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_1_comar1_G4_mul2_G16_mul1_G256_inv0 = (r00_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p1_0_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul1_G256_inv0);
    assign p0_G4_mul2_G16_mul1_G256_inv0 = (p0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign p1_G4_mul2_G16_mul1_G256_inv0 = (p1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul1_G256_inv0 = (r00_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r10_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r20_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r30_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r40_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul1_G256_inv0 = (r50_G4_mul2_G16_mul1_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul1_G256_inv0 = (b0_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul1_G256_inv0 = (d1_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul1_G256_inv0 = (d0_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign m3_comar2_G4_mul2_G16_mul1_G256_inv0 = (b1_G4_mul2_G16_mul1_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign p2_comar2_G4_mul2_G16_mul1_G256_inv0 = (m0_comar2_G4_mul2_G16_mul1_G256_inv0 & m1_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign p3_comar2_G4_mul2_G16_mul1_G256_inv0 = (m3_comar2_G4_mul2_G16_mul1_G256_inv0 & m2_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign p1_comar2_G4_mul2_G16_mul1_G256_inv0 = (m0_comar2_G4_mul2_G16_mul1_G256_inv0 & m2_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign p4_comar2_G4_mul2_G16_mul1_G256_inv0 = (m3_comar2_G4_mul2_G16_mul1_G256_inv0 & m1_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i0_comar2_G4_mul2_G16_mul1_G256_inv0 = (p1_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i1_comar2_G4_mul2_G16_mul1_G256_inv0 = (p2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i2_comar2_G4_mul2_G16_mul1_G256_inv0 = (p3_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i3_comar2_G4_mul2_G16_mul1_G256_inv0 = (p4_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0 = (i1_comar2_G4_mul2_G16_mul1_G256_inv0 ^ i2_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0 = (i0_comar2_G4_mul2_G16_mul1_G256_inv0 ^ i3_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign q0_0_G4_mul2_G16_mul1_G256_inv0 = (i1xori2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_1_comar2_G4_mul2_G16_mul1_G256_inv0 = (r00_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul1_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G4_mul2_G16_mul1_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul1_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G4_mul2_G16_mul1_G256_inv0 = (q0_0_G4_mul2_G16_mul1_G256_inv0 ^ e0_G4_mul2_G16_mul1_G256_inv0);
    assign q1_G4_mul2_G16_mul1_G256_inv0 = (q1_0_G4_mul2_G16_mul1_G256_inv0 ^ e1_G4_mul2_G16_mul1_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul1_G256_inv0 = (p1_G4_mul2_G16_mul1_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul2_G16_mul1_G256_inv0 = (p0_G4_mul2_G16_mul1_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul1_G256_inv0 = (p1ls1_G4_mul2_G16_mul1_G256_inv0 | q1_G4_mul2_G16_mul1_G256_inv0);
    assign q1_0_G16_mul1_G256_inv0 = (p0ls1_G4_mul2_G16_mul1_G256_inv0 | q0_G4_mul2_G16_mul1_G256_inv0);
    assign q0_G16_mul1_G256_inv0 = (q0_0_G16_mul1_G256_inv0 ^ e01_G16_mul1_G256_inv0);
    assign q1_G16_mul1_G256_inv0 = (q1_0_G16_mul1_G256_inv0 ^ e11_G16_mul1_G256_inv0);
    assign p0ls2_G16_mul1_G256_inv0 = (p0_G16_mul1_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_mul1_G256_inv0 = (p1_G16_mul1_G256_inv0 << dec_2_inp);
    assign p0_G256_inv0 = (p0ls2_G16_mul1_G256_inv0 | q0_G16_mul1_G256_inv0);
    assign p1_G256_inv0 = (p1ls2_G16_mul1_G256_inv0 | q1_G16_mul1_G256_inv0);
    assign r00_G16_mul2_G256_inv0 = (r0_inp % dec_16_inp);
    assign r10_G16_mul2_G256_inv0 = (r1_inp % dec_16_inp);
    assign r20_G16_mul2_G256_inv0 = (r2_inp % dec_16_inp);
    assign r30_G16_mul2_G256_inv0 = (r3_inp % dec_16_inp);
    assign r40_G16_mul2_G256_inv0 = (r4_inp % dec_16_inp);
    assign r50_G16_mul2_G256_inv0 = (r5_inp % dec_16_inp);
    assign a0_0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_12_inp);
    assign a1_0_G16_mul2_G256_inv0 = (e1_G256_inv0 & dec_12_inp);
    assign a0_G16_mul2_G256_inv0 = (a0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign a1_G16_mul2_G256_inv0 = (a1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign b0_G16_mul2_G256_inv0 = (e0_G256_inv0 & dec_3_inp);
    assign b1_G16_mul2_G256_inv0 = (e1_G256_inv0 & dec_3_inp);
    assign c0_0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_12_inp);
    assign c1_0_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_12_inp);
    assign c0_G16_mul2_G256_inv0 = (c0_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign c1_G16_mul2_G256_inv0 = (c1_0_G16_mul2_G256_inv0 >> dec_2_inp);
    assign d0_G16_mul2_G256_inv0 = (a0_G256_inv0 & dec_3_inp);
    assign d1_G16_mul2_G256_inv0 = (a1_G256_inv0 & dec_3_inp);
    assign axorb_0_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 ^ b0_G16_mul2_G256_inv0);
    assign cxord_0_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 ^ d0_G16_mul2_G256_inv0);
    assign axorb_1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 ^ b1_G16_mul2_G256_inv0);
    assign cxord_1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 ^ d1_G16_mul2_G256_inv0);
    assign r00_G4_mul0_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul0_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul0_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul0_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul0_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul0_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul0_G16_mul2_G256_inv0 = (a0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul0_G16_mul2_G256_inv0 = (a1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign b1_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul0_G16_mul2_G256_inv0 = (c0_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul0_G16_mul2_G256_inv0 = (c1_0_G4_mul0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ b0_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ d0_G4_mul0_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ b1_G4_mul0_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ d1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul0_G16_mul2_G256_inv0 = (axorb_0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul0_G16_mul2_G256_inv0 = (cxord_1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul0_G16_mul2_G256_inv0 = (cxord_0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign m3_comar0_G4_mul0_G16_mul2_G256_inv0 = (axorb_1_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign p2_comar0_G4_mul0_G16_mul2_G256_inv0 = (m0_comar0_G4_mul0_G16_mul2_G256_inv0 & m1_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign p3_comar0_G4_mul0_G16_mul2_G256_inv0 = (m3_comar0_G4_mul0_G16_mul2_G256_inv0 & m2_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_comar0_G4_mul0_G16_mul2_G256_inv0 = (m0_comar0_G4_mul0_G16_mul2_G256_inv0 & m2_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign p4_comar0_G4_mul0_G16_mul2_G256_inv0 = (m3_comar0_G4_mul0_G16_mul2_G256_inv0 & m1_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i0_comar0_G4_mul0_G16_mul2_G256_inv0 = (p1_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i1_comar0_G4_mul0_G16_mul2_G256_inv0 = (p2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i2_comar0_G4_mul0_G16_mul2_G256_inv0 = (p3_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i3_comar0_G4_mul0_G16_mul2_G256_inv0 = (p4_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0 = (i1_comar0_G4_mul0_G16_mul2_G256_inv0 ^ i2_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0 = (i0_comar0_G4_mul0_G16_mul2_G256_inv0 ^ i3_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign e0_G4_mul0_G16_mul2_G256_inv0 = (i1xori2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_1_comar0_G4_mul0_G16_mul2_G256_inv0 = (r00_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul0_G16_mul2_G256_inv0 = (a0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul0_G16_mul2_G256_inv0 = (c1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul0_G16_mul2_G256_inv0 = (c0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign m3_comar1_G4_mul0_G16_mul2_G256_inv0 = (a1_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p2_comar1_G4_mul0_G16_mul2_G256_inv0 = (m0_comar1_G4_mul0_G16_mul2_G256_inv0 & m1_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p3_comar1_G4_mul0_G16_mul2_G256_inv0 = (m3_comar1_G4_mul0_G16_mul2_G256_inv0 & m2_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p1_comar1_G4_mul0_G16_mul2_G256_inv0 = (m0_comar1_G4_mul0_G16_mul2_G256_inv0 & m2_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p4_comar1_G4_mul0_G16_mul2_G256_inv0 = (m3_comar1_G4_mul0_G16_mul2_G256_inv0 & m1_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i0_comar1_G4_mul0_G16_mul2_G256_inv0 = (p1_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i1_comar1_G4_mul0_G16_mul2_G256_inv0 = (p2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i2_comar1_G4_mul0_G16_mul2_G256_inv0 = (p3_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i3_comar1_G4_mul0_G16_mul2_G256_inv0 = (p4_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0 = (i1_comar1_G4_mul0_G16_mul2_G256_inv0 ^ i2_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0 = (i0_comar1_G4_mul0_G16_mul2_G256_inv0 ^ i3_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p0_0_G4_mul0_G16_mul2_G256_inv0 = (i1xori2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_1_comar1_G4_mul0_G16_mul2_G256_inv0 = (r00_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p1_0_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul0_G16_mul2_G256_inv0);
    assign p0_G4_mul0_G16_mul2_G256_inv0 = (p0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign p1_G4_mul0_G16_mul2_G256_inv0 = (p1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul0_G16_mul2_G256_inv0 = (r00_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r10_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r20_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r30_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r40_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul0_G16_mul2_G256_inv0 = (r50_G4_mul0_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul0_G16_mul2_G256_inv0 = (b0_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul0_G16_mul2_G256_inv0 = (d1_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul0_G16_mul2_G256_inv0 = (d0_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign m3_comar2_G4_mul0_G16_mul2_G256_inv0 = (b1_G4_mul0_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign p2_comar2_G4_mul0_G16_mul2_G256_inv0 = (m0_comar2_G4_mul0_G16_mul2_G256_inv0 & m1_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign p3_comar2_G4_mul0_G16_mul2_G256_inv0 = (m3_comar2_G4_mul0_G16_mul2_G256_inv0 & m2_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign p1_comar2_G4_mul0_G16_mul2_G256_inv0 = (m0_comar2_G4_mul0_G16_mul2_G256_inv0 & m2_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign p4_comar2_G4_mul0_G16_mul2_G256_inv0 = (m3_comar2_G4_mul0_G16_mul2_G256_inv0 & m1_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i0_comar2_G4_mul0_G16_mul2_G256_inv0 = (p1_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i1_comar2_G4_mul0_G16_mul2_G256_inv0 = (p2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i2_comar2_G4_mul0_G16_mul2_G256_inv0 = (p3_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i3_comar2_G4_mul0_G16_mul2_G256_inv0 = (p4_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0 = (i1_comar2_G4_mul0_G16_mul2_G256_inv0 ^ i2_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0 = (i0_comar2_G4_mul0_G16_mul2_G256_inv0 ^ i3_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign q0_0_G4_mul0_G16_mul2_G256_inv0 = (i1xori2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_1_comar2_G4_mul0_G16_mul2_G256_inv0 = (r00_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul0_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign q1_0_G4_mul0_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul0_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul0_G16_mul2_G256_inv0);
    assign q0_G4_mul0_G16_mul2_G256_inv0 = (q0_0_G4_mul0_G16_mul2_G256_inv0 ^ e0_G4_mul0_G16_mul2_G256_inv0);
    assign q1_G4_mul0_G16_mul2_G256_inv0 = (q1_0_G4_mul0_G16_mul2_G256_inv0 ^ e1_G4_mul0_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul0_G16_mul2_G256_inv0 = (p1_G4_mul0_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul0_G16_mul2_G256_inv0 = (p0_G4_mul0_G16_mul2_G256_inv0 << dec_1_inp);
    assign e0_G16_mul2_G256_inv0 = (p1ls1_G4_mul0_G16_mul2_G256_inv0 | q1_G4_mul0_G16_mul2_G256_inv0);
    assign e1_G16_mul2_G256_inv0 = (p0ls1_G4_mul0_G16_mul2_G256_inv0 | q0_G4_mul0_G16_mul2_G256_inv0);
    assign a0_0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a1_0_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_0_G4_scl_N0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign a1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_0_G4_scl_N0_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_scl_N0_G16_mul2_G256_inv0 = (e0_G16_mul2_G256_inv0 & dec_1_inp);
    assign b1_G4_scl_N0_G16_mul2_G256_inv0 = (e1_G16_mul2_G256_inv0 & dec_1_inp);
    assign p0_G4_scl_N0_G16_mul2_G256_inv0 = b0_G4_scl_N0_G16_mul2_G256_inv0;
    assign p1_G4_scl_N0_G16_mul2_G256_inv0 = b1_G4_scl_N0_G16_mul2_G256_inv0;
    assign q0_G4_scl_N0_G16_mul2_G256_inv0 = (a0_G4_scl_N0_G16_mul2_G256_inv0 ^ b0_G4_scl_N0_G16_mul2_G256_inv0);
    assign q1_G4_scl_N0_G16_mul2_G256_inv0 = (a1_G4_scl_N0_G16_mul2_G256_inv0 ^ b1_G4_scl_N0_G16_mul2_G256_inv0);
    assign p1ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p1_G4_scl_N0_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_scl_N0_G16_mul2_G256_inv0 = (p0_G4_scl_N0_G16_mul2_G256_inv0 << dec_1_inp);
    assign e01_G16_mul2_G256_inv0 = (p0ls1_G4_scl_N0_G16_mul2_G256_inv0 | q0_G4_scl_N0_G16_mul2_G256_inv0);
    assign e11_G16_mul2_G256_inv0 = (p1ls1_G4_scl_N0_G16_mul2_G256_inv0 | q1_G4_scl_N0_G16_mul2_G256_inv0);
    assign r00_G4_mul1_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul1_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul1_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul1_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul1_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul1_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul1_G16_mul2_G256_inv0 = (a0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul1_G16_mul2_G256_inv0 = (a1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul1_G16_mul2_G256_inv0 = (a0_G16_mul2_G256_inv0 & dec_1_inp);
    assign b1_G4_mul1_G16_mul2_G256_inv0 = (a1_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul1_G16_mul2_G256_inv0 = (c0_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul1_G16_mul2_G256_inv0 = (c1_0_G4_mul1_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul1_G16_mul2_G256_inv0 = (c0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul1_G16_mul2_G256_inv0 = (c1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ b0_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ d0_G4_mul1_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ b1_G4_mul1_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ d1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul1_G16_mul2_G256_inv0 = (axorb_0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul1_G16_mul2_G256_inv0 = (cxord_1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul1_G16_mul2_G256_inv0 = (cxord_0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign m3_comar0_G4_mul1_G16_mul2_G256_inv0 = (axorb_1_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign p2_comar0_G4_mul1_G16_mul2_G256_inv0 = (m0_comar0_G4_mul1_G16_mul2_G256_inv0 & m1_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign p3_comar0_G4_mul1_G16_mul2_G256_inv0 = (m3_comar0_G4_mul1_G16_mul2_G256_inv0 & m2_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_comar0_G4_mul1_G16_mul2_G256_inv0 = (m0_comar0_G4_mul1_G16_mul2_G256_inv0 & m2_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign p4_comar0_G4_mul1_G16_mul2_G256_inv0 = (m3_comar0_G4_mul1_G16_mul2_G256_inv0 & m1_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i0_comar0_G4_mul1_G16_mul2_G256_inv0 = (p1_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i1_comar0_G4_mul1_G16_mul2_G256_inv0 = (p2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i2_comar0_G4_mul1_G16_mul2_G256_inv0 = (p3_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i3_comar0_G4_mul1_G16_mul2_G256_inv0 = (p4_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0 = (i1_comar0_G4_mul1_G16_mul2_G256_inv0 ^ i2_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0 = (i0_comar0_G4_mul1_G16_mul2_G256_inv0 ^ i3_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign e0_G4_mul1_G16_mul2_G256_inv0 = (i1xori2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_1_comar0_G4_mul1_G16_mul2_G256_inv0 = (r00_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign e1_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul1_G16_mul2_G256_inv0 = (a0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul1_G16_mul2_G256_inv0 = (c1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul1_G16_mul2_G256_inv0 = (c0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign m3_comar1_G4_mul1_G16_mul2_G256_inv0 = (a1_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p2_comar1_G4_mul1_G16_mul2_G256_inv0 = (m0_comar1_G4_mul1_G16_mul2_G256_inv0 & m1_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p3_comar1_G4_mul1_G16_mul2_G256_inv0 = (m3_comar1_G4_mul1_G16_mul2_G256_inv0 & m2_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_comar1_G4_mul1_G16_mul2_G256_inv0 = (m0_comar1_G4_mul1_G16_mul2_G256_inv0 & m2_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p4_comar1_G4_mul1_G16_mul2_G256_inv0 = (m3_comar1_G4_mul1_G16_mul2_G256_inv0 & m1_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i0_comar1_G4_mul1_G16_mul2_G256_inv0 = (p1_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i1_comar1_G4_mul1_G16_mul2_G256_inv0 = (p2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i2_comar1_G4_mul1_G16_mul2_G256_inv0 = (p3_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i3_comar1_G4_mul1_G16_mul2_G256_inv0 = (p4_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0 = (i1_comar1_G4_mul1_G16_mul2_G256_inv0 ^ i2_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0 = (i0_comar1_G4_mul1_G16_mul2_G256_inv0 ^ i3_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p0_0_G4_mul1_G16_mul2_G256_inv0 = (i1xori2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_1_comar1_G4_mul1_G16_mul2_G256_inv0 = (r00_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G4_mul1_G16_mul2_G256_inv0 = (p0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign p1_G4_mul1_G16_mul2_G256_inv0 = (p1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul1_G16_mul2_G256_inv0 = (r00_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r10_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r20_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r30_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r40_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul1_G16_mul2_G256_inv0 = (r50_G4_mul1_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul1_G16_mul2_G256_inv0 = (b0_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul1_G16_mul2_G256_inv0 = (d1_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul1_G16_mul2_G256_inv0 = (d0_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign m3_comar2_G4_mul1_G16_mul2_G256_inv0 = (b1_G4_mul1_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign p2_comar2_G4_mul1_G16_mul2_G256_inv0 = (m0_comar2_G4_mul1_G16_mul2_G256_inv0 & m1_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign p3_comar2_G4_mul1_G16_mul2_G256_inv0 = (m3_comar2_G4_mul1_G16_mul2_G256_inv0 & m2_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign p1_comar2_G4_mul1_G16_mul2_G256_inv0 = (m0_comar2_G4_mul1_G16_mul2_G256_inv0 & m2_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign p4_comar2_G4_mul1_G16_mul2_G256_inv0 = (m3_comar2_G4_mul1_G16_mul2_G256_inv0 & m1_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i0_comar2_G4_mul1_G16_mul2_G256_inv0 = (p1_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i1_comar2_G4_mul1_G16_mul2_G256_inv0 = (p2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i2_comar2_G4_mul1_G16_mul2_G256_inv0 = (p3_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i3_comar2_G4_mul1_G16_mul2_G256_inv0 = (p4_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0 = (i1_comar2_G4_mul1_G16_mul2_G256_inv0 ^ i2_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0 = (i0_comar2_G4_mul1_G16_mul2_G256_inv0 ^ i3_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign q0_0_G4_mul1_G16_mul2_G256_inv0 = (i1xori2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_1_comar2_G4_mul1_G16_mul2_G256_inv0 = (r00_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul1_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign q1_0_G4_mul1_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul1_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul1_G16_mul2_G256_inv0);
    assign q0_G4_mul1_G16_mul2_G256_inv0 = (q0_0_G4_mul1_G16_mul2_G256_inv0 ^ e0_G4_mul1_G16_mul2_G256_inv0);
    assign q1_G4_mul1_G16_mul2_G256_inv0 = (q1_0_G4_mul1_G16_mul2_G256_inv0 ^ e1_G4_mul1_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul1_G16_mul2_G256_inv0 = (p1_G4_mul1_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul1_G16_mul2_G256_inv0 = (p0_G4_mul1_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul1_G16_mul2_G256_inv0 | q1_G4_mul1_G16_mul2_G256_inv0);
    assign p1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul1_G16_mul2_G256_inv0 | q0_G4_mul1_G16_mul2_G256_inv0);
    assign p0_G16_mul2_G256_inv0 = (p0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign p1_G16_mul2_G256_inv0 = (p1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign r00_G4_mul2_G16_mul2_G256_inv0 = (r00_G16_mul2_G256_inv0 % dec_4_inp);
    assign r10_G4_mul2_G16_mul2_G256_inv0 = (r10_G16_mul2_G256_inv0 % dec_4_inp);
    assign r20_G4_mul2_G16_mul2_G256_inv0 = (r20_G16_mul2_G256_inv0 % dec_4_inp);
    assign r30_G4_mul2_G16_mul2_G256_inv0 = (r30_G16_mul2_G256_inv0 % dec_4_inp);
    assign r40_G4_mul2_G16_mul2_G256_inv0 = (r40_G16_mul2_G256_inv0 % dec_4_inp);
    assign r50_G4_mul2_G16_mul2_G256_inv0 = (r50_G16_mul2_G256_inv0 % dec_4_inp);
    assign a0_0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_2_inp);
    assign a1_0_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & dec_2_inp);
    assign a0_G4_mul2_G16_mul2_G256_inv0 = (a0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign a1_G4_mul2_G16_mul2_G256_inv0 = (a1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign b0_G4_mul2_G16_mul2_G256_inv0 = (b0_G16_mul2_G256_inv0 & dec_1_inp);
    assign b1_G4_mul2_G16_mul2_G256_inv0 = (b1_G16_mul2_G256_inv0 & dec_1_inp);
    assign c0_0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_2_inp);
    assign c1_0_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_2_inp);
    assign c0_G4_mul2_G16_mul2_G256_inv0 = (c0_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign c1_G4_mul2_G16_mul2_G256_inv0 = (c1_0_G4_mul2_G16_mul2_G256_inv0 >> dec_1_inp);
    assign d0_G4_mul2_G16_mul2_G256_inv0 = (d0_G16_mul2_G256_inv0 & dec_1_inp);
    assign d1_G4_mul2_G16_mul2_G256_inv0 = (d1_G16_mul2_G256_inv0 & dec_1_inp);
    assign axorb_0_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ b0_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_0_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ d0_G4_mul2_G16_mul2_G256_inv0);
    assign axorb_1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ b1_G4_mul2_G16_mul2_G256_inv0);
    assign cxord_1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ d1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar0_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar0_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar0_G4_mul2_G16_mul2_G256_inv0 = (axorb_0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar0_G4_mul2_G16_mul2_G256_inv0 = (cxord_1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar0_G4_mul2_G16_mul2_G256_inv0 = (cxord_0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign m3_comar0_G4_mul2_G16_mul2_G256_inv0 = (axorb_1_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign p2_comar0_G4_mul2_G16_mul2_G256_inv0 = (m0_comar0_G4_mul2_G16_mul2_G256_inv0 & m1_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign p3_comar0_G4_mul2_G16_mul2_G256_inv0 = (m3_comar0_G4_mul2_G16_mul2_G256_inv0 & m2_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_comar0_G4_mul2_G16_mul2_G256_inv0 = (m0_comar0_G4_mul2_G16_mul2_G256_inv0 & m2_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign p4_comar0_G4_mul2_G16_mul2_G256_inv0 = (m3_comar0_G4_mul2_G16_mul2_G256_inv0 & m1_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i0_comar0_G4_mul2_G16_mul2_G256_inv0 = (p1_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i1_comar0_G4_mul2_G16_mul2_G256_inv0 = (p2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i2_comar0_G4_mul2_G16_mul2_G256_inv0 = (p3_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i3_comar0_G4_mul2_G16_mul2_G256_inv0 = (p4_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0 = (i1_comar0_G4_mul2_G16_mul2_G256_inv0 ^ i2_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0 = (i0_comar0_G4_mul2_G16_mul2_G256_inv0 ^ i3_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign e0_G4_mul2_G16_mul2_G256_inv0 = (i1xori2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_1_comar0_G4_mul2_G16_mul2_G256_inv0 = (r00_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar0_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign e1_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar0_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar0_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar1_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar1_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar1_G4_mul2_G16_mul2_G256_inv0 = (a0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar1_G4_mul2_G16_mul2_G256_inv0 = (c1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar1_G4_mul2_G16_mul2_G256_inv0 = (c0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign m3_comar1_G4_mul2_G16_mul2_G256_inv0 = (a1_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p2_comar1_G4_mul2_G16_mul2_G256_inv0 = (m0_comar1_G4_mul2_G16_mul2_G256_inv0 & m1_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p3_comar1_G4_mul2_G16_mul2_G256_inv0 = (m3_comar1_G4_mul2_G16_mul2_G256_inv0 & m2_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p1_comar1_G4_mul2_G16_mul2_G256_inv0 = (m0_comar1_G4_mul2_G16_mul2_G256_inv0 & m2_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p4_comar1_G4_mul2_G16_mul2_G256_inv0 = (m3_comar1_G4_mul2_G16_mul2_G256_inv0 & m1_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i0_comar1_G4_mul2_G16_mul2_G256_inv0 = (p1_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i1_comar1_G4_mul2_G16_mul2_G256_inv0 = (p2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i2_comar1_G4_mul2_G16_mul2_G256_inv0 = (p3_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i3_comar1_G4_mul2_G16_mul2_G256_inv0 = (p4_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0 = (i1_comar1_G4_mul2_G16_mul2_G256_inv0 ^ i2_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0 = (i0_comar1_G4_mul2_G16_mul2_G256_inv0 ^ i3_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p0_0_G4_mul2_G16_mul2_G256_inv0 = (i1xori2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_1_comar1_G4_mul2_G16_mul2_G256_inv0 = (r00_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar1_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p1_0_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar1_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar1_G4_mul2_G16_mul2_G256_inv0);
    assign p0_G4_mul2_G16_mul2_G256_inv0 = (p0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign p1_G4_mul2_G16_mul2_G256_inv0 = (p1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign r00_comar2_G4_mul2_G16_mul2_G256_inv0 = (r00_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r10_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r0_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r20_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r1_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r30_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r2_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r40_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign r3_10_comar2_G4_mul2_G16_mul2_G256_inv0 = (r50_G4_mul2_G16_mul2_G256_inv0 % dec_2_inp);
    assign m0_comar2_G4_mul2_G16_mul2_G256_inv0 = (b0_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign m1_comar2_G4_mul2_G16_mul2_G256_inv0 = (d1_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign m2_comar2_G4_mul2_G16_mul2_G256_inv0 = (d0_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign m3_comar2_G4_mul2_G16_mul2_G256_inv0 = (b1_G4_mul2_G16_mul2_G256_inv0 ^ r00_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign p2_comar2_G4_mul2_G16_mul2_G256_inv0 = (m0_comar2_G4_mul2_G16_mul2_G256_inv0 & m1_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign p3_comar2_G4_mul2_G16_mul2_G256_inv0 = (m3_comar2_G4_mul2_G16_mul2_G256_inv0 & m2_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign p1_comar2_G4_mul2_G16_mul2_G256_inv0 = (m0_comar2_G4_mul2_G16_mul2_G256_inv0 & m2_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign p4_comar2_G4_mul2_G16_mul2_G256_inv0 = (m3_comar2_G4_mul2_G16_mul2_G256_inv0 & m1_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i0_comar2_G4_mul2_G16_mul2_G256_inv0 = (p1_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i1_comar2_G4_mul2_G16_mul2_G256_inv0 = (p2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i2_comar2_G4_mul2_G16_mul2_G256_inv0 = (p3_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i3_comar2_G4_mul2_G16_mul2_G256_inv0 = (p4_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0 = (i1_comar2_G4_mul2_G16_mul2_G256_inv0 ^ i2_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0 = (i0_comar2_G4_mul2_G16_mul2_G256_inv0 ^ i3_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign q0_0_G4_mul2_G16_mul2_G256_inv0 = (i1xori2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ i0xori3_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_1_comar2_G4_mul2_G16_mul2_G256_inv0 = (r00_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_2_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_1_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r0_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_3_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_2_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r1_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign y1_4_comar2_G4_mul2_G16_mul2_G256_inv0 = (y1_3_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r2_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G4_mul2_G16_mul2_G256_inv0 = (y1_4_comar2_G4_mul2_G16_mul2_G256_inv0 ^ r3_10_comar2_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G4_mul2_G16_mul2_G256_inv0 = (q0_0_G4_mul2_G16_mul2_G256_inv0 ^ e0_G4_mul2_G16_mul2_G256_inv0);
    assign q1_G4_mul2_G16_mul2_G256_inv0 = (q1_0_G4_mul2_G16_mul2_G256_inv0 ^ e1_G4_mul2_G16_mul2_G256_inv0);
    assign p1ls1_G4_mul2_G16_mul2_G256_inv0 = (p1_G4_mul2_G16_mul2_G256_inv0 << dec_1_inp);
    assign p0ls1_G4_mul2_G16_mul2_G256_inv0 = (p0_G4_mul2_G16_mul2_G256_inv0 << dec_1_inp);
    assign q0_0_G16_mul2_G256_inv0 = (p1ls1_G4_mul2_G16_mul2_G256_inv0 | q1_G4_mul2_G16_mul2_G256_inv0);
    assign q1_0_G16_mul2_G256_inv0 = (p0ls1_G4_mul2_G16_mul2_G256_inv0 | q0_G4_mul2_G16_mul2_G256_inv0);
    assign q0_G16_mul2_G256_inv0 = (q0_0_G16_mul2_G256_inv0 ^ e01_G16_mul2_G256_inv0);
    assign q1_G16_mul2_G256_inv0 = (q1_0_G16_mul2_G256_inv0 ^ e11_G16_mul2_G256_inv0);
    assign p0ls2_G16_mul2_G256_inv0 = (p0_G16_mul2_G256_inv0 << dec_2_inp);
    assign p1ls2_G16_mul2_G256_inv0 = (p1_G16_mul2_G256_inv0 << dec_2_inp);
    assign q0_G256_inv0 = (p0ls2_G16_mul2_G256_inv0 | q0_G16_mul2_G256_inv0);
    assign q1_G256_inv0 = (p1ls2_G16_mul2_G256_inv0 | q1_G16_mul2_G256_inv0);
    assign p0ls4_G256_inv0 = (p0_G256_inv0 << dec_4_inp);
    assign p1ls4_G256_inv0 = (p1_G256_inv0 << dec_4_inp);
    assign t4 = (p0ls4_G256_inv0 | q0_G256_inv0);
    assign t5 = (p1ls4_G256_inv0 | q1_G256_inv0);
    assign y_G256_newbasis1 = dec_0_inp;
    assign tempy1_G256_newbasis1 = y_G256_newbasis1;
    assign cond1_G256_newbasis1 = (t4 & dec_1_inp);
    assign negCond1_G256_newbasis1 = !cond1_G256_newbasis1;
    assign yxorb1_G256_newbasis1 = (y_G256_newbasis1 ^ dec_36_inp);
    assign ny1_G256_newbasis1 = (cond1_G256_newbasis1 * yxorb1_G256_newbasis1);
    assign tempybooloNegCond1_G256_newbasis1 = (tempy1_G256_newbasis1 * negCond1_G256_newbasis1);
    assign y1_G256_newbasis1 = (ny1_G256_newbasis1 + tempybooloNegCond1_G256_newbasis1);
    assign x1_G256_newbasis1 = (t4 >> dec_1_inp);
    assign tempy2_G256_newbasis1 = y1_G256_newbasis1;
    assign cond2_G256_newbasis1 = (x1_G256_newbasis1 & dec_1_inp);
    assign negCond2_G256_newbasis1 = !cond2_G256_newbasis1;
    assign yxorb2_G256_newbasis1 = (y1_G256_newbasis1 ^ dec_3_inp);
    assign ny2_G256_newbasis1 = (cond2_G256_newbasis1 * yxorb2_G256_newbasis1);
    assign tempybooloNegCond2_G256_newbasis1 = (tempy2_G256_newbasis1 * negCond2_G256_newbasis1);
    assign y2_G256_newbasis1 = (ny2_G256_newbasis1 + tempybooloNegCond2_G256_newbasis1);
    assign x2_G256_newbasis1 = (x1_G256_newbasis1 >> dec_1_inp);
    assign tempy3_G256_newbasis1 = y2_G256_newbasis1;
    assign cond3_G256_newbasis1 = (x2_G256_newbasis1 & dec_1_inp);
    assign negCond3_G256_newbasis1 = !cond3_G256_newbasis1;
    assign yxorb3_G256_newbasis1 = (y2_G256_newbasis1 ^ dec_4_inp);
    assign ny3_G256_newbasis1 = (cond3_G256_newbasis1 * yxorb3_G256_newbasis1);
    assign tempybooloNegCond3_G256_newbasis1 = (tempy3_G256_newbasis1 * negCond3_G256_newbasis1);
    assign y3_G256_newbasis1 = (ny3_G256_newbasis1 + tempybooloNegCond3_G256_newbasis1);
    assign x3_G256_newbasis1 = (x2_G256_newbasis1 >> dec_1_inp);
    assign tempy4_G256_newbasis1 = y3_G256_newbasis1;
    assign cond4_G256_newbasis1 = (x3_G256_newbasis1 & dec_1_inp);
    assign negCond4_G256_newbasis1 = !cond4_G256_newbasis1;
    assign yxorb4_G256_newbasis1 = (y3_G256_newbasis1 ^ dec_220_inp);
    assign ny4_G256_newbasis1 = (cond4_G256_newbasis1 * yxorb4_G256_newbasis1);
    assign tempybooloNegCond4_G256_newbasis1 = (tempy4_G256_newbasis1 * negCond4_G256_newbasis1);
    assign y4_G256_newbasis1 = (ny4_G256_newbasis1 + tempybooloNegCond4_G256_newbasis1);
    assign x4_G256_newbasis1 = (x3_G256_newbasis1 >> dec_1_inp);
    assign tempy5_G256_newbasis1 = y4_G256_newbasis1;
    assign cond5_G256_newbasis1 = (x4_G256_newbasis1 & dec_1_inp);
    assign negCond5_G256_newbasis1 = !cond5_G256_newbasis1;
    assign yxorb5_G256_newbasis1 = (y4_G256_newbasis1 ^ dec_11_inp);
    assign ny5_G256_newbasis1 = (cond5_G256_newbasis1 * yxorb5_G256_newbasis1);
    assign tempybooloNegCond5_G256_newbasis1 = (tempy5_G256_newbasis1 * negCond5_G256_newbasis1);
    assign y5_G256_newbasis1 = (ny5_G256_newbasis1 + tempybooloNegCond5_G256_newbasis1);
    assign x5_G256_newbasis1 = (x4_G256_newbasis1 >> dec_1_inp);
    assign tempy6_G256_newbasis1 = y5_G256_newbasis1;
    assign cond6_G256_newbasis1 = (x5_G256_newbasis1 & dec_1_inp);
    assign negCond6_G256_newbasis1 = !cond6_G256_newbasis1;
    assign yxorb6_G256_newbasis1 = (y5_G256_newbasis1 ^ dec_158_inp);
    assign ny6_G256_newbasis1 = (cond6_G256_newbasis1 * yxorb6_G256_newbasis1);
    assign tempybooloNegCond6_G256_newbasis1 = (tempy6_G256_newbasis1 * negCond6_G256_newbasis1);
    assign y6_G256_newbasis1 = (ny6_G256_newbasis1 + tempybooloNegCond6_G256_newbasis1);
    assign x6_G256_newbasis1 = (x5_G256_newbasis1 >> dec_1_inp);
    assign tempy7_G256_newbasis1 = y6_G256_newbasis1;
    assign cond7_G256_newbasis1 = (x6_G256_newbasis1 & dec_1_inp);
    assign negCond7_G256_newbasis1 = !cond7_G256_newbasis1;
    assign yxorb7_G256_newbasis1 = (y6_G256_newbasis1 ^ dec_45_inp);
    assign ny7_G256_newbasis1 = (cond7_G256_newbasis1 * yxorb7_G256_newbasis1);
    assign tempybooloNegCond7_G256_newbasis1 = (tempy7_G256_newbasis1 * negCond7_G256_newbasis1);
    assign y7_G256_newbasis1 = (ny7_G256_newbasis1 + tempybooloNegCond7_G256_newbasis1);
    assign x7_G256_newbasis1 = (x6_G256_newbasis1 >> dec_1_inp);
    assign tempy8_G256_newbasis1 = y7_G256_newbasis1;
    assign cond8_G256_newbasis1 = (x7_G256_newbasis1 & dec_1_inp);
    assign negCond8_G256_newbasis1 = !cond8_G256_newbasis1;
    assign yxorb8_G256_newbasis1 = (y7_G256_newbasis1 ^ dec_88_inp);
    assign ny8_G256_newbasis1 = (cond8_G256_newbasis1 * yxorb8_G256_newbasis1);
    assign tempybooloNegCond8_G256_newbasis1 = (tempy8_G256_newbasis1 * negCond8_G256_newbasis1);
    assign y8_G256_newbasis1 = (ny8_G256_newbasis1 + tempybooloNegCond8_G256_newbasis1);
    assign x8_G256_newbasis1 = (x7_G256_newbasis1 >> dec_1_inp);
    assign t6 = y8_G256_newbasis1;
    assign z_y_G256_newbasis1 = dec_0_inp;
    assign z_tempy1_G256_newbasis1 = z_y_G256_newbasis1;
    assign z_cond1_G256_newbasis1 = (t5 & dec_1_inp);
    assign z_negCond1_G256_newbasis1 = !z_cond1_G256_newbasis1;
    assign z_yxorb1_G256_newbasis1 = (z_y_G256_newbasis1 ^ dec_36_inp);
    assign z_ny1_G256_newbasis1 = (z_cond1_G256_newbasis1 * z_yxorb1_G256_newbasis1);
    assign z_tempybooloNegCond1_G256_newbasis1 = (z_tempy1_G256_newbasis1 * z_negCond1_G256_newbasis1);
    assign z_y1_G256_newbasis1 = (z_ny1_G256_newbasis1 + z_tempybooloNegCond1_G256_newbasis1);
    assign z_x1_G256_newbasis1 = (t5 >> dec_1_inp);
    assign z_tempy2_G256_newbasis1 = z_y1_G256_newbasis1;
    assign z_cond2_G256_newbasis1 = (z_x1_G256_newbasis1 & dec_1_inp);
    assign z_negCond2_G256_newbasis1 = !z_cond2_G256_newbasis1;
    assign z_yxorb2_G256_newbasis1 = (z_y1_G256_newbasis1 ^ dec_3_inp);
    assign z_ny2_G256_newbasis1 = (z_cond2_G256_newbasis1 * z_yxorb2_G256_newbasis1);
    assign z_tempybooloNegCond2_G256_newbasis1 = (z_tempy2_G256_newbasis1 * z_negCond2_G256_newbasis1);
    assign z_y2_G256_newbasis1 = (z_ny2_G256_newbasis1 + z_tempybooloNegCond2_G256_newbasis1);
    assign z_x2_G256_newbasis1 = (z_x1_G256_newbasis1 >> dec_1_inp);
    assign z_tempy3_G256_newbasis1 = z_y2_G256_newbasis1;
    assign z_cond3_G256_newbasis1 = (z_x2_G256_newbasis1 & dec_1_inp);
    assign z_negCond3_G256_newbasis1 = !z_cond3_G256_newbasis1;
    assign z_yxorb3_G256_newbasis1 = (z_y2_G256_newbasis1 ^ dec_4_inp);
    assign z_ny3_G256_newbasis1 = (z_cond3_G256_newbasis1 * z_yxorb3_G256_newbasis1);
    assign z_tempybooloNegCond3_G256_newbasis1 = (z_tempy3_G256_newbasis1 * z_negCond3_G256_newbasis1);
    assign z_y3_G256_newbasis1 = (z_ny3_G256_newbasis1 + z_tempybooloNegCond3_G256_newbasis1);
    assign z_x3_G256_newbasis1 = (z_x2_G256_newbasis1 >> dec_1_inp);
    assign z_tempy4_G256_newbasis1 = z_y3_G256_newbasis1;
    assign z_cond4_G256_newbasis1 = (z_x3_G256_newbasis1 & dec_1_inp);
    assign z_negCond4_G256_newbasis1 = !z_cond4_G256_newbasis1;
    assign z_yxorb4_G256_newbasis1 = (z_y3_G256_newbasis1 ^ dec_220_inp);
    assign z_ny4_G256_newbasis1 = (z_cond4_G256_newbasis1 * z_yxorb4_G256_newbasis1);
    assign z_tempybooloNegCond4_G256_newbasis1 = (z_tempy4_G256_newbasis1 * z_negCond4_G256_newbasis1);
    assign z_y4_G256_newbasis1 = (z_ny4_G256_newbasis1 + z_tempybooloNegCond4_G256_newbasis1);
    assign z_x4_G256_newbasis1 = (z_x3_G256_newbasis1 >> dec_1_inp);
    assign z_tempy5_G256_newbasis1 = z_y4_G256_newbasis1;
    assign z_cond5_G256_newbasis1 = (z_x4_G256_newbasis1 & dec_1_inp);
    assign z_negCond5_G256_newbasis1 = !z_cond5_G256_newbasis1;
    assign z_yxorb5_G256_newbasis1 = (z_y4_G256_newbasis1 ^ dec_11_inp);
    assign z_ny5_G256_newbasis1 = (z_cond5_G256_newbasis1 * z_yxorb5_G256_newbasis1);
    assign z_tempybooloNegCond5_G256_newbasis1 = (z_tempy5_G256_newbasis1 * z_negCond5_G256_newbasis1);
    assign z_y5_G256_newbasis1 = (z_ny5_G256_newbasis1 + z_tempybooloNegCond5_G256_newbasis1);
    assign z_x5_G256_newbasis1 = (z_x4_G256_newbasis1 >> dec_1_inp);
    assign z_tempy6_G256_newbasis1 = z_y5_G256_newbasis1;
    assign z_cond6_G256_newbasis1 = (z_x5_G256_newbasis1 & dec_1_inp);
    assign z_negCond6_G256_newbasis1 = !z_cond6_G256_newbasis1;
    assign z_yxorb6_G256_newbasis1 = (z_y5_G256_newbasis1 ^ dec_158_inp);
    assign z_ny6_G256_newbasis1 = (z_cond6_G256_newbasis1 * z_yxorb6_G256_newbasis1);
    assign z_tempybooloNegCond6_G256_newbasis1 = (z_tempy6_G256_newbasis1 * z_negCond6_G256_newbasis1);
    assign z_y6_G256_newbasis1 = (z_ny6_G256_newbasis1 + z_tempybooloNegCond6_G256_newbasis1);
    assign z_x6_G256_newbasis1 = (z_x5_G256_newbasis1 >> dec_1_inp);
    assign z_tempy7_G256_newbasis1 = z_y6_G256_newbasis1;
    assign z_cond7_G256_newbasis1 = (z_x6_G256_newbasis1 & dec_1_inp);
    assign z_negCond7_G256_newbasis1 = !z_cond7_G256_newbasis1;
    assign z_yxorb7_G256_newbasis1 = (z_y6_G256_newbasis1 ^ dec_45_inp);
    assign z_ny7_G256_newbasis1 = (z_cond7_G256_newbasis1 * z_yxorb7_G256_newbasis1);
    assign z_tempybooloNegCond7_G256_newbasis1 = (z_tempy7_G256_newbasis1 * z_negCond7_G256_newbasis1);
    assign z_y7_G256_newbasis1 = (z_ny7_G256_newbasis1 + z_tempybooloNegCond7_G256_newbasis1);
    assign z_x7_G256_newbasis1 = (z_x6_G256_newbasis1 >> dec_1_inp);
    assign z_tempy8_G256_newbasis1 = z_y7_G256_newbasis1;
    assign z_cond8_G256_newbasis1 = (z_x7_G256_newbasis1 & dec_1_inp);
    assign z_negCond8_G256_newbasis1 = !z_cond8_G256_newbasis1;
    assign z_yxorb8_G256_newbasis1 = (z_y7_G256_newbasis1 ^ dec_88_inp);
    assign z_ny8_G256_newbasis1 = (z_cond8_G256_newbasis1 * z_yxorb8_G256_newbasis1);
    assign z_tempybooloNegCond8_G256_newbasis1 = (z_tempy8_G256_newbasis1 * z_negCond8_G256_newbasis1);
    assign z_y8_G256_newbasis1 = (z_ny8_G256_newbasis1 + z_tempybooloNegCond8_G256_newbasis1);
    assign z_x8_G256_newbasis1 = (z_x7_G256_newbasis1 >> dec_1_inp);
    assign t7 = z_y8_G256_newbasis1;

    always @(posedge clk) begin
        y0 <= (t6 ^ dec_99_inp);
        y1 <= t7;
    end

endmodule

